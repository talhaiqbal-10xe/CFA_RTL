`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:49:42 08/03/2022 
// Design Name: 
// Module Name:    equ_24_27_comp 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: This module needs equ_24_27 as well as pre_equ_24_27
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module equ_24_27_comp(
    );


endmodule
