module adder4x19(
output [20:0] out1,out2,
input [18:0]A,B,C,D );


wire [21:0] CV;
 assign CV=21'b000000000000000000010;




///////////// Iteration Number =1///////////////////





wire Hi1L0_inp1, Hi1L0_inp2;
assign Hi1L0_inp1 = A[0];
assign Hi1L0_inp2 = B[0];
wire sHi1L0, cHi1L0;
HA Hi1L0 ( sHi1L0,cHi1L0,Hi1L0_inp1,Hi1L0_inp2 );

wire F1i1L1_inp1, F1i1L1_inp2, F1i1L1_inp3;
assign F1i1L1_inp1 = A[1];
assign F1i1L1_inp2 = B[1];
assign F1i1L1_inp3 = C[1];
wire sF1i1L1, cF1i1L1;
FA F1i1L1( sF1i1L1,cF1i1L1,F1i1L1_inp1,F1i1L1_inp2,F1i1L1_inp3 );

wire Hi1L1_inp1, Hi1L1_inp2;
assign Hi1L1_inp1 = D[1];
assign Hi1L1_inp2 = CV[1];
wire sHi1L1, cHi1L1;
HA Hi1L1 ( sHi1L1,cHi1L1,Hi1L1_inp1,Hi1L1_inp2 );

wire F1i1L2_inp1, F1i1L2_inp2, F1i1L2_inp3;
assign F1i1L2_inp1 = A[2];
assign F1i1L2_inp2 = B[2];
assign F1i1L2_inp3 = C[2];
wire sF1i1L2, cF1i1L2;
FA F1i1L2( sF1i1L2,cF1i1L2,F1i1L2_inp1,F1i1L2_inp2,F1i1L2_inp3 );

wire Hi1L2_inp1, Hi1L2_inp2;
assign Hi1L2_inp1 = D[2];
assign Hi1L2_inp2 = cF1i1L1;
wire sHi1L2, cHi1L2;
HA Hi1L2 ( sHi1L2,cHi1L2,Hi1L2_inp1,Hi1L2_inp2 );

wire F1i1L3_inp1, F1i1L3_inp2, F1i1L3_inp3;
assign F1i1L3_inp1 = A[3];
assign F1i1L3_inp2 = B[3];
assign F1i1L3_inp3 = C[3];
wire sF1i1L3, cF1i1L3;
FA F1i1L3( sF1i1L3,cF1i1L3,F1i1L3_inp1,F1i1L3_inp2,F1i1L3_inp3 );

wire Hi1L3_inp1, Hi1L3_inp2;
assign Hi1L3_inp1 = D[3];
assign Hi1L3_inp2 = cF1i1L2;
wire sHi1L3, cHi1L3;
HA Hi1L3 ( sHi1L3,cHi1L3,Hi1L3_inp1,Hi1L3_inp2 );

wire F1i1L4_inp1, F1i1L4_inp2, F1i1L4_inp3;
assign F1i1L4_inp1 = A[4];
assign F1i1L4_inp2 = B[4];
assign F1i1L4_inp3 = C[4];
wire sF1i1L4, cF1i1L4;
FA F1i1L4( sF1i1L4,cF1i1L4,F1i1L4_inp1,F1i1L4_inp2,F1i1L4_inp3 );

wire Hi1L4_inp1, Hi1L4_inp2;
assign Hi1L4_inp1 = D[4];
assign Hi1L4_inp2 = cF1i1L3;
wire sHi1L4, cHi1L4;
HA Hi1L4 ( sHi1L4,cHi1L4,Hi1L4_inp1,Hi1L4_inp2 );

wire F1i1L5_inp1, F1i1L5_inp2, F1i1L5_inp3;
assign F1i1L5_inp1 = A[5];
assign F1i1L5_inp2 = B[5];
assign F1i1L5_inp3 = C[5];
wire sF1i1L5, cF1i1L5;
FA F1i1L5( sF1i1L5,cF1i1L5,F1i1L5_inp1,F1i1L5_inp2,F1i1L5_inp3 );

wire Hi1L5_inp1, Hi1L5_inp2;
assign Hi1L5_inp1 = D[5];
assign Hi1L5_inp2 = cF1i1L4;
wire sHi1L5, cHi1L5;
HA Hi1L5 ( sHi1L5,cHi1L5,Hi1L5_inp1,Hi1L5_inp2 );

wire F1i1L6_inp1, F1i1L6_inp2, F1i1L6_inp3;
assign F1i1L6_inp1 = A[6];
assign F1i1L6_inp2 = B[6];
assign F1i1L6_inp3 = C[6];
wire sF1i1L6, cF1i1L6;
FA F1i1L6( sF1i1L6,cF1i1L6,F1i1L6_inp1,F1i1L6_inp2,F1i1L6_inp3 );

wire Hi1L6_inp1, Hi1L6_inp2;
assign Hi1L6_inp1 = D[6];
assign Hi1L6_inp2 = cF1i1L5;
wire sHi1L6, cHi1L6;
HA Hi1L6 ( sHi1L6,cHi1L6,Hi1L6_inp1,Hi1L6_inp2 );

wire F1i1L7_inp1, F1i1L7_inp2, F1i1L7_inp3;
assign F1i1L7_inp1 = A[7];
assign F1i1L7_inp2 = B[7];
assign F1i1L7_inp3 = C[7];
wire sF1i1L7, cF1i1L7;
FA F1i1L7( sF1i1L7,cF1i1L7,F1i1L7_inp1,F1i1L7_inp2,F1i1L7_inp3 );

wire Hi1L7_inp1, Hi1L7_inp2;
assign Hi1L7_inp1 = D[7];
assign Hi1L7_inp2 = cF1i1L6;
wire sHi1L7, cHi1L7;
HA Hi1L7 ( sHi1L7,cHi1L7,Hi1L7_inp1,Hi1L7_inp2 );

wire F1i1L8_inp1, F1i1L8_inp2, F1i1L8_inp3;
assign F1i1L8_inp1 = A[8];
assign F1i1L8_inp2 = B[8];
assign F1i1L8_inp3 = C[8];
wire sF1i1L8, cF1i1L8;
FA F1i1L8( sF1i1L8,cF1i1L8,F1i1L8_inp1,F1i1L8_inp2,F1i1L8_inp3 );

wire Hi1L8_inp1, Hi1L8_inp2;
assign Hi1L8_inp1 = D[8];
assign Hi1L8_inp2 = cF1i1L7;
wire sHi1L8, cHi1L8;
HA Hi1L8 ( sHi1L8,cHi1L8,Hi1L8_inp1,Hi1L8_inp2 );

wire F1i1L9_inp1, F1i1L9_inp2, F1i1L9_inp3;
assign F1i1L9_inp1 = A[9];
assign F1i1L9_inp2 = B[9];
assign F1i1L9_inp3 = C[9];
wire sF1i1L9, cF1i1L9;
FA F1i1L9( sF1i1L9,cF1i1L9,F1i1L9_inp1,F1i1L9_inp2,F1i1L9_inp3 );

wire Hi1L9_inp1, Hi1L9_inp2;
assign Hi1L9_inp1 = D[9];
assign Hi1L9_inp2 = cF1i1L8;
wire sHi1L9, cHi1L9;
HA Hi1L9 ( sHi1L9,cHi1L9,Hi1L9_inp1,Hi1L9_inp2 );

wire F1i1L10_inp1, F1i1L10_inp2, F1i1L10_inp3;
assign F1i1L10_inp1 = A[10];
assign F1i1L10_inp2 = B[10];
assign F1i1L10_inp3 = C[10];
wire sF1i1L10, cF1i1L10;
FA F1i1L10( sF1i1L10,cF1i1L10,F1i1L10_inp1,F1i1L10_inp2,F1i1L10_inp3 );

wire Hi1L10_inp1, Hi1L10_inp2;
assign Hi1L10_inp1 = D[10];
assign Hi1L10_inp2 = cF1i1L9;
wire sHi1L10, cHi1L10;
HA Hi1L10 ( sHi1L10,cHi1L10,Hi1L10_inp1,Hi1L10_inp2 );

wire F1i1L11_inp1, F1i1L11_inp2, F1i1L11_inp3;
assign F1i1L11_inp1 = A[11];
assign F1i1L11_inp2 = B[11];
assign F1i1L11_inp3 = C[11];
wire sF1i1L11, cF1i1L11;
FA F1i1L11( sF1i1L11,cF1i1L11,F1i1L11_inp1,F1i1L11_inp2,F1i1L11_inp3 );

wire Hi1L11_inp1, Hi1L11_inp2;
assign Hi1L11_inp1 = D[11];
assign Hi1L11_inp2 = cF1i1L10;
wire sHi1L11, cHi1L11;
HA Hi1L11 ( sHi1L11,cHi1L11,Hi1L11_inp1,Hi1L11_inp2 );

wire F1i1L12_inp1, F1i1L12_inp2, F1i1L12_inp3;
assign F1i1L12_inp1 = A[12];
assign F1i1L12_inp2 = B[12];
assign F1i1L12_inp3 = C[12];
wire sF1i1L12, cF1i1L12;
FA F1i1L12( sF1i1L12,cF1i1L12,F1i1L12_inp1,F1i1L12_inp2,F1i1L12_inp3 );

wire Hi1L12_inp1, Hi1L12_inp2;
assign Hi1L12_inp1 = D[12];
assign Hi1L12_inp2 = cF1i1L11;
wire sHi1L12, cHi1L12;
HA Hi1L12 ( sHi1L12,cHi1L12,Hi1L12_inp1,Hi1L12_inp2 );

wire F1i1L13_inp1, F1i1L13_inp2, F1i1L13_inp3;
assign F1i1L13_inp1 = A[13];
assign F1i1L13_inp2 = B[13];
assign F1i1L13_inp3 = C[13];
wire sF1i1L13, cF1i1L13;
FA F1i1L13( sF1i1L13,cF1i1L13,F1i1L13_inp1,F1i1L13_inp2,F1i1L13_inp3 );

wire Hi1L13_inp1, Hi1L13_inp2;
assign Hi1L13_inp1 = D[13];
assign Hi1L13_inp2 = cF1i1L12;
wire sHi1L13, cHi1L13;
HA Hi1L13 ( sHi1L13,cHi1L13,Hi1L13_inp1,Hi1L13_inp2 );

wire F1i1L14_inp1, F1i1L14_inp2, F1i1L14_inp3;
assign F1i1L14_inp1 = A[14];
assign F1i1L14_inp2 = B[14];
assign F1i1L14_inp3 = C[14];
wire sF1i1L14, cF1i1L14;
FA F1i1L14( sF1i1L14,cF1i1L14,F1i1L14_inp1,F1i1L14_inp2,F1i1L14_inp3 );

wire Hi1L14_inp1, Hi1L14_inp2;
assign Hi1L14_inp1 = D[14];
assign Hi1L14_inp2 = cF1i1L13;
wire sHi1L14, cHi1L14;
HA Hi1L14 ( sHi1L14,cHi1L14,Hi1L14_inp1,Hi1L14_inp2 );

wire F1i1L15_inp1, F1i1L15_inp2, F1i1L15_inp3;
assign F1i1L15_inp1 = A[15];
assign F1i1L15_inp2 = B[15];
assign F1i1L15_inp3 = C[15];
wire sF1i1L15, cF1i1L15;
FA F1i1L15( sF1i1L15,cF1i1L15,F1i1L15_inp1,F1i1L15_inp2,F1i1L15_inp3 );

wire Hi1L15_inp1, Hi1L15_inp2;
assign Hi1L15_inp1 = D[15];
assign Hi1L15_inp2 = cF1i1L14;
wire sHi1L15, cHi1L15;
HA Hi1L15 ( sHi1L15,cHi1L15,Hi1L15_inp1,Hi1L15_inp2 );

wire F1i1L16_inp1, F1i1L16_inp2, F1i1L16_inp3;
assign F1i1L16_inp1 = A[16];
assign F1i1L16_inp2 = B[16];
assign F1i1L16_inp3 = C[16];
wire sF1i1L16, cF1i1L16;
FA F1i1L16( sF1i1L16,cF1i1L16,F1i1L16_inp1,F1i1L16_inp2,F1i1L16_inp3 );

wire Hi1L16_inp1, Hi1L16_inp2;
assign Hi1L16_inp1 = D[16];
assign Hi1L16_inp2 = cF1i1L15;
wire sHi1L16, cHi1L16;
HA Hi1L16 ( sHi1L16,cHi1L16,Hi1L16_inp1,Hi1L16_inp2 );

wire F1i1L17_inp1, F1i1L17_inp2, F1i1L17_inp3;
assign F1i1L17_inp1 = A[17];
assign F1i1L17_inp2 = B[17];
assign F1i1L17_inp3 = C[17];
wire sF1i1L17, cF1i1L17;
FA F1i1L17( sF1i1L17,cF1i1L17,F1i1L17_inp1,F1i1L17_inp2,F1i1L17_inp3 );

wire Hi1L17_inp1, Hi1L17_inp2;
assign Hi1L17_inp1 = D[17];
assign Hi1L17_inp2 = cF1i1L16;
wire sHi1L17, cHi1L17;
HA Hi1L17 ( sHi1L17,cHi1L17,Hi1L17_inp1,Hi1L17_inp2 );

wire F1i1L18_inp1, F1i1L18_inp2, F1i1L18_inp3;
assign F1i1L18_inp1 = A[18];
assign F1i1L18_inp2 = B[18];
assign F1i1L18_inp3 = C[18];
wire sF1i1L18, cF1i1L18;
FA F1i1L18( sF1i1L18,cF1i1L18,F1i1L18_inp1,F1i1L18_inp2,F1i1L18_inp3 );

wire Hi1L18_inp1, Hi1L18_inp2;
assign Hi1L18_inp1 = D[18];
assign Hi1L18_inp2 = cF1i1L17;
wire sHi1L18, cHi1L18;
HA Hi1L18 ( sHi1L18,cHi1L18,Hi1L18_inp1,Hi1L18_inp2 );



///////////// Iteration Number =2///////////////////





wire Hi2L0_inp1, Hi2L0_inp2;
assign Hi2L0_inp1 = C[0];
assign Hi2L0_inp2 = D[0];
wire sHi2L0, cHi2L0;
HA Hi2L0 ( sHi2L0,cHi2L0,Hi2L0_inp1,Hi2L0_inp2 );

wire F1i2L1_inp1, F1i2L1_inp2, F1i2L1_inp3;
assign F1i2L1_inp1 = cHi1L0;
assign F1i2L1_inp2 = sF1i1L1;
assign F1i2L1_inp3 = sHi1L1;
wire sF1i2L1, cF1i2L1;
FA F1i2L1( sF1i2L1,cF1i2L1,F1i2L1_inp1,F1i2L1_inp2,F1i2L1_inp3 );

wire F1i2L2_inp1, F1i2L2_inp2, F1i2L2_inp3;
assign F1i2L2_inp1 = cHi1L1;
assign F1i2L2_inp2 = sF1i1L2;
assign F1i2L2_inp3 = sHi1L2;
wire sF1i2L2, cF1i2L2;
FA F1i2L2( sF1i2L2,cF1i2L2,F1i2L2_inp1,F1i2L2_inp2,F1i2L2_inp3 );

wire F1i2L3_inp1, F1i2L3_inp2, F1i2L3_inp3;
assign F1i2L3_inp1 = cHi1L2;
assign F1i2L3_inp2 = sF1i1L3;
assign F1i2L3_inp3 = sHi1L3;
wire sF1i2L3, cF1i2L3;
FA F1i2L3( sF1i2L3,cF1i2L3,F1i2L3_inp1,F1i2L3_inp2,F1i2L3_inp3 );

wire F1i2L4_inp1, F1i2L4_inp2, F1i2L4_inp3;
assign F1i2L4_inp1 = cHi1L3;
assign F1i2L4_inp2 = sF1i1L4;
assign F1i2L4_inp3 = sHi1L4;
wire sF1i2L4, cF1i2L4;
FA F1i2L4( sF1i2L4,cF1i2L4,F1i2L4_inp1,F1i2L4_inp2,F1i2L4_inp3 );

wire F1i2L5_inp1, F1i2L5_inp2, F1i2L5_inp3;
assign F1i2L5_inp1 = cHi1L4;
assign F1i2L5_inp2 = sF1i1L5;
assign F1i2L5_inp3 = sHi1L5;
wire sF1i2L5, cF1i2L5;
FA F1i2L5( sF1i2L5,cF1i2L5,F1i2L5_inp1,F1i2L5_inp2,F1i2L5_inp3 );

wire F1i2L6_inp1, F1i2L6_inp2, F1i2L6_inp3;
assign F1i2L6_inp1 = cHi1L5;
assign F1i2L6_inp2 = sF1i1L6;
assign F1i2L6_inp3 = sHi1L6;
wire sF1i2L6, cF1i2L6;
FA F1i2L6( sF1i2L6,cF1i2L6,F1i2L6_inp1,F1i2L6_inp2,F1i2L6_inp3 );

wire F1i2L7_inp1, F1i2L7_inp2, F1i2L7_inp3;
assign F1i2L7_inp1 = cHi1L6;
assign F1i2L7_inp2 = sF1i1L7;
assign F1i2L7_inp3 = sHi1L7;
wire sF1i2L7, cF1i2L7;
FA F1i2L7( sF1i2L7,cF1i2L7,F1i2L7_inp1,F1i2L7_inp2,F1i2L7_inp3 );

wire F1i2L8_inp1, F1i2L8_inp2, F1i2L8_inp3;
assign F1i2L8_inp1 = cHi1L7;
assign F1i2L8_inp2 = sF1i1L8;
assign F1i2L8_inp3 = sHi1L8;
wire sF1i2L8, cF1i2L8;
FA F1i2L8( sF1i2L8,cF1i2L8,F1i2L8_inp1,F1i2L8_inp2,F1i2L8_inp3 );

wire F1i2L9_inp1, F1i2L9_inp2, F1i2L9_inp3;
assign F1i2L9_inp1 = cHi1L8;
assign F1i2L9_inp2 = sF1i1L9;
assign F1i2L9_inp3 = sHi1L9;
wire sF1i2L9, cF1i2L9;
FA F1i2L9( sF1i2L9,cF1i2L9,F1i2L9_inp1,F1i2L9_inp2,F1i2L9_inp3 );

wire F1i2L10_inp1, F1i2L10_inp2, F1i2L10_inp3;
assign F1i2L10_inp1 = cHi1L9;
assign F1i2L10_inp2 = sF1i1L10;
assign F1i2L10_inp3 = sHi1L10;
wire sF1i2L10, cF1i2L10;
FA F1i2L10( sF1i2L10,cF1i2L10,F1i2L10_inp1,F1i2L10_inp2,F1i2L10_inp3 );

wire F1i2L11_inp1, F1i2L11_inp2, F1i2L11_inp3;
assign F1i2L11_inp1 = cHi1L10;
assign F1i2L11_inp2 = sF1i1L11;
assign F1i2L11_inp3 = sHi1L11;
wire sF1i2L11, cF1i2L11;
FA F1i2L11( sF1i2L11,cF1i2L11,F1i2L11_inp1,F1i2L11_inp2,F1i2L11_inp3 );

wire F1i2L12_inp1, F1i2L12_inp2, F1i2L12_inp3;
assign F1i2L12_inp1 = cHi1L11;
assign F1i2L12_inp2 = sF1i1L12;
assign F1i2L12_inp3 = sHi1L12;
wire sF1i2L12, cF1i2L12;
FA F1i2L12( sF1i2L12,cF1i2L12,F1i2L12_inp1,F1i2L12_inp2,F1i2L12_inp3 );

wire F1i2L13_inp1, F1i2L13_inp2, F1i2L13_inp3;
assign F1i2L13_inp1 = cHi1L12;
assign F1i2L13_inp2 = sF1i1L13;
assign F1i2L13_inp3 = sHi1L13;
wire sF1i2L13, cF1i2L13;
FA F1i2L13( sF1i2L13,cF1i2L13,F1i2L13_inp1,F1i2L13_inp2,F1i2L13_inp3 );

wire F1i2L14_inp1, F1i2L14_inp2, F1i2L14_inp3;
assign F1i2L14_inp1 = cHi1L13;
assign F1i2L14_inp2 = sF1i1L14;
assign F1i2L14_inp3 = sHi1L14;
wire sF1i2L14, cF1i2L14;
FA F1i2L14( sF1i2L14,cF1i2L14,F1i2L14_inp1,F1i2L14_inp2,F1i2L14_inp3 );

wire F1i2L15_inp1, F1i2L15_inp2, F1i2L15_inp3;
assign F1i2L15_inp1 = cHi1L14;
assign F1i2L15_inp2 = sF1i1L15;
assign F1i2L15_inp3 = sHi1L15;
wire sF1i2L15, cF1i2L15;
FA F1i2L15( sF1i2L15,cF1i2L15,F1i2L15_inp1,F1i2L15_inp2,F1i2L15_inp3 );

wire F1i2L16_inp1, F1i2L16_inp2, F1i2L16_inp3;
assign F1i2L16_inp1 = cHi1L15;
assign F1i2L16_inp2 = sF1i1L16;
assign F1i2L16_inp3 = sHi1L16;
wire sF1i2L16, cF1i2L16;
FA F1i2L16( sF1i2L16,cF1i2L16,F1i2L16_inp1,F1i2L16_inp2,F1i2L16_inp3 );

wire F1i2L17_inp1, F1i2L17_inp2, F1i2L17_inp3;
assign F1i2L17_inp1 = cHi1L16;
assign F1i2L17_inp2 = sF1i1L17;
assign F1i2L17_inp3 = sHi1L17;
wire sF1i2L17, cF1i2L17;
FA F1i2L17( sF1i2L17,cF1i2L17,F1i2L17_inp1,F1i2L17_inp2,F1i2L17_inp3 );

wire F1i2L18_inp1, F1i2L18_inp2, F1i2L18_inp3;
assign F1i2L18_inp1 = cHi1L17;
assign F1i2L18_inp2 = sF1i1L18;
assign F1i2L18_inp3 = sHi1L18;
wire sF1i2L18, cF1i2L18;
FA F1i2L18( sF1i2L18,cF1i2L18,F1i2L18_inp1,F1i2L18_inp2,F1i2L18_inp3 );

wire Hi2L19_inp1, Hi2L19_inp2;
assign Hi2L19_inp1 = cF1i1L18;
assign Hi2L19_inp2 = cHi1L18;
wire sHi2L19, cHi2L19;
HA Hi2L19 ( sHi2L19,cHi2L19,Hi2L19_inp1,Hi2L19_inp2 );


assign out1 ={{cHi2L19},{cF1i2L18},{cF1i2L17},{cF1i2L16},{cF1i2L15},{cF1i2L14},{cF1i2L13},{cF1i2L12},{cF1i2L11},{cF1i2L10},{cF1i2L9},{cF1i2L8},{cF1i2L7},{cF1i2L6},{cF1i2L5},{cF1i2L4},{cF1i2L3},{cF1i2L2},{cF1i2L1},{cHi2L0},{sHi1L0}};
assign out2 ={{1'b0},{sHi2L19},{sF1i2L18},{sF1i2L17},{sF1i2L16},{sF1i2L15},{sF1i2L14},{sF1i2L13},{sF1i2L12},{sF1i2L11},{sF1i2L10},{sF1i2L9},{sF1i2L8},{sF1i2L7},{sF1i2L6},{sF1i2L5},{sF1i2L4},{sF1i2L3},{sF1i2L2},{sF1i2L1},{sHi2L0}} ;
endmodule