module mult11x11MAC(
output [21:0] out1,out2,
input [10:0] A,
input [10:0] B,
input [10:0]C );


integer i;
 reg[10:0] PP[ 0:10];
always@*
begin
   for ( i=0 ; i<11; i = i+1 )
   begin
      PP[i]= A & {11{B[i]}};
   end
end



///////////// Iteration Number =1///////////////////





wire Hi1L8_inp1, Hi1L8_inp2;
assign Hi1L8_inp1 = PP[0][8];
assign Hi1L8_inp2 = PP[1][7];
wire sHi1L8, cHi1L8;
HA Hi1L8 ( sHi1L8,cHi1L8,Hi1L8_inp1,Hi1L8_inp2 );

wire F1i1L9_inp1, F1i1L9_inp2, F1i1L9_inp3;
assign F1i1L9_inp1 = PP[0][9];
assign F1i1L9_inp2 = PP[1][8];
assign F1i1L9_inp3 = PP[2][7];
wire sF1i1L9, cF1i1L9;
FA F1i1L9( sF1i1L9,cF1i1L9,F1i1L9_inp1,F1i1L9_inp2,F1i1L9_inp3 );

wire Hi1L9_inp1, Hi1L9_inp2;
assign Hi1L9_inp1 = PP[3][6];
assign Hi1L9_inp2 = PP[4][5];
wire sHi1L9, cHi1L9;
HA Hi1L9 ( sHi1L9,cHi1L9,Hi1L9_inp1,Hi1L9_inp2 );

wire F1i1L10_inp1, F1i1L10_inp2, F1i1L10_inp3;
assign F1i1L10_inp1 = PP[0][10];
assign F1i1L10_inp2 = PP[1][9];
assign F1i1L10_inp3 = PP[2][8];
wire sF1i1L10, cF1i1L10;
FA F1i1L10( sF1i1L10,cF1i1L10,F1i1L10_inp1,F1i1L10_inp2,F1i1L10_inp3 );

wire F2i1L10_inp1, F2i1L10_inp2, F2i1L10_inp3;
assign F2i1L10_inp1 = PP[3][7];
assign F2i1L10_inp2 = PP[4][6];
assign F2i1L10_inp3 = PP[5][5];
wire sF2i1L10, cF2i1L10;
FA F2i1L10( sF2i1L10,cF2i1L10,F2i1L10_inp1,F2i1L10_inp2,F2i1L10_inp3 );

wire Hi1L10_inp1, Hi1L10_inp2;
assign Hi1L10_inp1 = PP[6][4];
assign Hi1L10_inp2 = PP[7][3];
wire sHi1L10, cHi1L10;
HA Hi1L10 ( sHi1L10,cHi1L10,Hi1L10_inp1,Hi1L10_inp2 );

wire F1i1L11_inp1, F1i1L11_inp2, F1i1L11_inp3;
assign F1i1L11_inp1 = PP[1][10];
assign F1i1L11_inp2 = PP[2][9];
assign F1i1L11_inp3 = PP[3][8];
wire sF1i1L11, cF1i1L11;
FA F1i1L11( sF1i1L11,cF1i1L11,F1i1L11_inp1,F1i1L11_inp2,F1i1L11_inp3 );

wire F2i1L11_inp1, F2i1L11_inp2, F2i1L11_inp3;
assign F2i1L11_inp1 = PP[4][7];
assign F2i1L11_inp2 = PP[5][6];
assign F2i1L11_inp3 = PP[6][5];
wire sF2i1L11, cF2i1L11;
FA F2i1L11( sF2i1L11,cF2i1L11,F2i1L11_inp1,F2i1L11_inp2,F2i1L11_inp3 );

wire F1i1L12_inp1, F1i1L12_inp2, F1i1L12_inp3;
assign F1i1L12_inp1 = PP[2][10];
assign F1i1L12_inp2 = PP[3][9];
assign F1i1L12_inp3 = PP[4][8];
wire sF1i1L12, cF1i1L12;
FA F1i1L12( sF1i1L12,cF1i1L12,F1i1L12_inp1,F1i1L12_inp2,F1i1L12_inp3 );



///////////// Iteration Number =2///////////////////





wire Hi2L5_inp1, Hi2L5_inp2;
assign Hi2L5_inp1 = PP[0][5];
assign Hi2L5_inp2 = PP[1][4];
wire sHi2L5, cHi2L5;
HA Hi2L5 ( sHi2L5,cHi2L5,Hi2L5_inp1,Hi2L5_inp2 );

wire F1i2L6_inp1, F1i2L6_inp2, F1i2L6_inp3;
assign F1i2L6_inp1 = PP[0][6];
assign F1i2L6_inp2 = PP[1][5];
assign F1i2L6_inp3 = PP[2][4];
wire sF1i2L6, cF1i2L6;
FA F1i2L6( sF1i2L6,cF1i2L6,F1i2L6_inp1,F1i2L6_inp2,F1i2L6_inp3 );

wire Hi2L6_inp1, Hi2L6_inp2;
assign Hi2L6_inp1 = PP[3][3];
assign Hi2L6_inp2 = PP[4][2];
wire sHi2L6, cHi2L6;
HA Hi2L6 ( sHi2L6,cHi2L6,Hi2L6_inp1,Hi2L6_inp2 );

wire F1i2L7_inp1, F1i2L7_inp2, F1i2L7_inp3;
assign F1i2L7_inp1 = PP[0][7];
assign F1i2L7_inp2 = PP[1][6];
assign F1i2L7_inp3 = PP[2][5];
wire sF1i2L7, cF1i2L7;
FA F1i2L7( sF1i2L7,cF1i2L7,F1i2L7_inp1,F1i2L7_inp2,F1i2L7_inp3 );

wire F2i2L7_inp1, F2i2L7_inp2, F2i2L7_inp3;
assign F2i2L7_inp1 = PP[3][4];
assign F2i2L7_inp2 = PP[4][3];
assign F2i2L7_inp3 = PP[5][2];
wire sF2i2L7, cF2i2L7;
FA F2i2L7( sF2i2L7,cF2i2L7,F2i2L7_inp1,F2i2L7_inp2,F2i2L7_inp3 );

wire Hi2L7_inp1, Hi2L7_inp2;
assign Hi2L7_inp1 = PP[6][1];
assign Hi2L7_inp2 = PP[7][0];
wire sHi2L7, cHi2L7;
HA Hi2L7 ( sHi2L7,cHi2L7,Hi2L7_inp1,Hi2L7_inp2 );

wire F1i2L8_inp1, F1i2L8_inp2, F1i2L8_inp3;
assign F1i2L8_inp1 = PP[2][6];
assign F1i2L8_inp2 = PP[3][5];
assign F1i2L8_inp3 = PP[4][4];
wire sF1i2L8, cF1i2L8;
FA F1i2L8( sF1i2L8,cF1i2L8,F1i2L8_inp1,F1i2L8_inp2,F1i2L8_inp3 );

wire F2i2L8_inp1, F2i2L8_inp2, F2i2L8_inp3;
assign F2i2L8_inp1 = PP[5][3];
assign F2i2L8_inp2 = PP[6][2];
assign F2i2L8_inp3 = PP[7][1];
wire sF2i2L8, cF2i2L8;
FA F2i2L8( sF2i2L8,cF2i2L8,F2i2L8_inp1,F2i2L8_inp2,F2i2L8_inp3 );

wire F3i2L8_inp1, F3i2L8_inp2, F3i2L8_inp3;
assign F3i2L8_inp1 = PP[8][0];
assign F3i2L8_inp2 = C[8];
assign F3i2L8_inp3 = sHi1L8;
wire sF3i2L8, cF3i2L8;
FA F3i2L8( sF3i2L8,cF3i2L8,F3i2L8_inp1,F3i2L8_inp2,F3i2L8_inp3 );

wire F1i2L9_inp1, F1i2L9_inp2, F1i2L9_inp3;
assign F1i2L9_inp1 = PP[5][4];
assign F1i2L9_inp2 = PP[6][3];
assign F1i2L9_inp3 = PP[7][2];
wire sF1i2L9, cF1i2L9;
FA F1i2L9( sF1i2L9,cF1i2L9,F1i2L9_inp1,F1i2L9_inp2,F1i2L9_inp3 );

wire F2i2L9_inp1, F2i2L9_inp2, F2i2L9_inp3;
assign F2i2L9_inp1 = PP[8][1];
assign F2i2L9_inp2 = PP[9][0];
assign F2i2L9_inp3 = C[9];
wire sF2i2L9, cF2i2L9;
FA F2i2L9( sF2i2L9,cF2i2L9,F2i2L9_inp1,F2i2L9_inp2,F2i2L9_inp3 );

wire F3i2L9_inp1, F3i2L9_inp2, F3i2L9_inp3;
assign F3i2L9_inp1 = cHi1L8;
assign F3i2L9_inp2 = sF1i1L9;
assign F3i2L9_inp3 = sHi1L9;
wire sF3i2L9, cF3i2L9;
FA F3i2L9( sF3i2L9,cF3i2L9,F3i2L9_inp1,F3i2L9_inp2,F3i2L9_inp3 );

wire F1i2L10_inp1, F1i2L10_inp2, F1i2L10_inp3;
assign F1i2L10_inp1 = PP[8][2];
assign F1i2L10_inp2 = PP[9][1];
assign F1i2L10_inp3 = PP[10][0];
wire sF1i2L10, cF1i2L10;
FA F1i2L10( sF1i2L10,cF1i2L10,F1i2L10_inp1,F1i2L10_inp2,F1i2L10_inp3 );

wire F2i2L10_inp1, F2i2L10_inp2, F2i2L10_inp3;
assign F2i2L10_inp1 = C[10];
assign F2i2L10_inp2 = cF1i1L9;
assign F2i2L10_inp3 = cHi1L9;
wire sF2i2L10, cF2i2L10;
FA F2i2L10( sF2i2L10,cF2i2L10,F2i2L10_inp1,F2i2L10_inp2,F2i2L10_inp3 );

wire F3i2L10_inp1, F3i2L10_inp2, F3i2L10_inp3;
assign F3i2L10_inp1 = sF1i1L10;
assign F3i2L10_inp2 = sF2i1L10;
assign F3i2L10_inp3 = sHi1L10;
wire sF3i2L10, cF3i2L10;
FA F3i2L10( sF3i2L10,cF3i2L10,F3i2L10_inp1,F3i2L10_inp2,F3i2L10_inp3 );

wire F1i2L11_inp1, F1i2L11_inp2, F1i2L11_inp3;
assign F1i2L11_inp1 = PP[7][4];
assign F1i2L11_inp2 = PP[8][3];
assign F1i2L11_inp3 = PP[9][2];
wire sF1i2L11, cF1i2L11;
FA F1i2L11( sF1i2L11,cF1i2L11,F1i2L11_inp1,F1i2L11_inp2,F1i2L11_inp3 );

wire F2i2L11_inp1, F2i2L11_inp2, F2i2L11_inp3;
assign F2i2L11_inp1 = PP[10][1];
assign F2i2L11_inp2 = cF1i1L10;
assign F2i2L11_inp3 = cF2i1L10;
wire sF2i2L11, cF2i2L11;
FA F2i2L11( sF2i2L11,cF2i2L11,F2i2L11_inp1,F2i2L11_inp2,F2i2L11_inp3 );

wire F3i2L11_inp1, F3i2L11_inp2, F3i2L11_inp3;
assign F3i2L11_inp1 = cHi1L10;
assign F3i2L11_inp2 = sF1i1L11;
assign F3i2L11_inp3 = sF2i1L11;
wire sF3i2L11, cF3i2L11;
FA F3i2L11( sF3i2L11,cF3i2L11,F3i2L11_inp1,F3i2L11_inp2,F3i2L11_inp3 );

wire F1i2L12_inp1, F1i2L12_inp2, F1i2L12_inp3;
assign F1i2L12_inp1 = PP[5][7];
assign F1i2L12_inp2 = PP[6][6];
assign F1i2L12_inp3 = PP[7][5];
wire sF1i2L12, cF1i2L12;
FA F1i2L12( sF1i2L12,cF1i2L12,F1i2L12_inp1,F1i2L12_inp2,F1i2L12_inp3 );

wire F2i2L12_inp1, F2i2L12_inp2, F2i2L12_inp3;
assign F2i2L12_inp1 = PP[8][4];
assign F2i2L12_inp2 = PP[9][3];
assign F2i2L12_inp3 = PP[10][2];
wire sF2i2L12, cF2i2L12;
FA F2i2L12( sF2i2L12,cF2i2L12,F2i2L12_inp1,F2i2L12_inp2,F2i2L12_inp3 );

wire F3i2L12_inp1, F3i2L12_inp2, F3i2L12_inp3;
assign F3i2L12_inp1 = cF1i1L11;
assign F3i2L12_inp2 = cF2i1L11;
assign F3i2L12_inp3 = sF1i1L12;
wire sF3i2L12, cF3i2L12;
FA F3i2L12( sF3i2L12,cF3i2L12,F3i2L12_inp1,F3i2L12_inp2,F3i2L12_inp3 );

wire F1i2L13_inp1, F1i2L13_inp2, F1i2L13_inp3;
assign F1i2L13_inp1 = PP[3][10];
assign F1i2L13_inp2 = PP[4][9];
assign F1i2L13_inp3 = PP[5][8];
wire sF1i2L13, cF1i2L13;
FA F1i2L13( sF1i2L13,cF1i2L13,F1i2L13_inp1,F1i2L13_inp2,F1i2L13_inp3 );

wire F2i2L13_inp1, F2i2L13_inp2, F2i2L13_inp3;
assign F2i2L13_inp1 = PP[6][7];
assign F2i2L13_inp2 = PP[7][6];
assign F2i2L13_inp3 = PP[8][5];
wire sF2i2L13, cF2i2L13;
FA F2i2L13( sF2i2L13,cF2i2L13,F2i2L13_inp1,F2i2L13_inp2,F2i2L13_inp3 );

wire F3i2L13_inp1, F3i2L13_inp2, F3i2L13_inp3;
assign F3i2L13_inp1 = PP[9][4];
assign F3i2L13_inp2 = PP[10][3];
assign F3i2L13_inp3 = cF1i1L12;
wire sF3i2L13, cF3i2L13;
FA F3i2L13( sF3i2L13,cF3i2L13,F3i2L13_inp1,F3i2L13_inp2,F3i2L13_inp3 );

wire F1i2L14_inp1, F1i2L14_inp2, F1i2L14_inp3;
assign F1i2L14_inp1 = PP[4][10];
assign F1i2L14_inp2 = PP[5][9];
assign F1i2L14_inp3 = PP[6][8];
wire sF1i2L14, cF1i2L14;
FA F1i2L14( sF1i2L14,cF1i2L14,F1i2L14_inp1,F1i2L14_inp2,F1i2L14_inp3 );

wire F2i2L14_inp1, F2i2L14_inp2, F2i2L14_inp3;
assign F2i2L14_inp1 = PP[7][7];
assign F2i2L14_inp2 = PP[8][6];
assign F2i2L14_inp3 = PP[9][5];
wire sF2i2L14, cF2i2L14;
FA F2i2L14( sF2i2L14,cF2i2L14,F2i2L14_inp1,F2i2L14_inp2,F2i2L14_inp3 );

wire F1i2L15_inp1, F1i2L15_inp2, F1i2L15_inp3;
assign F1i2L15_inp1 = PP[5][10];
assign F1i2L15_inp2 = PP[6][9];
assign F1i2L15_inp3 = PP[7][8];
wire sF1i2L15, cF1i2L15;
FA F1i2L15( sF1i2L15,cF1i2L15,F1i2L15_inp1,F1i2L15_inp2,F1i2L15_inp3 );



///////////// Iteration Number =3///////////////////





wire Hi3L3_inp1, Hi3L3_inp2;
assign Hi3L3_inp1 = PP[0][3];
assign Hi3L3_inp2 = PP[1][2];
wire sHi3L3, cHi3L3;
HA Hi3L3 ( sHi3L3,cHi3L3,Hi3L3_inp1,Hi3L3_inp2 );

wire F1i3L4_inp1, F1i3L4_inp2, F1i3L4_inp3;
assign F1i3L4_inp1 = PP[0][4];
assign F1i3L4_inp2 = PP[1][3];
assign F1i3L4_inp3 = PP[2][2];
wire sF1i3L4, cF1i3L4;
FA F1i3L4( sF1i3L4,cF1i3L4,F1i3L4_inp1,F1i3L4_inp2,F1i3L4_inp3 );

wire Hi3L4_inp1, Hi3L4_inp2;
assign Hi3L4_inp1 = PP[3][1];
assign Hi3L4_inp2 = PP[4][0];
wire sHi3L4, cHi3L4;
HA Hi3L4 ( sHi3L4,cHi3L4,Hi3L4_inp1,Hi3L4_inp2 );

wire F1i3L5_inp1, F1i3L5_inp2, F1i3L5_inp3;
assign F1i3L5_inp1 = PP[2][3];
assign F1i3L5_inp2 = PP[3][2];
assign F1i3L5_inp3 = PP[4][1];
wire sF1i3L5, cF1i3L5;
FA F1i3L5( sF1i3L5,cF1i3L5,F1i3L5_inp1,F1i3L5_inp2,F1i3L5_inp3 );

wire F2i3L5_inp1, F2i3L5_inp2, F2i3L5_inp3;
assign F2i3L5_inp1 = PP[5][0];
assign F2i3L5_inp2 = C[5];
assign F2i3L5_inp3 = sHi2L5;
wire sF2i3L5, cF2i3L5;
FA F2i3L5( sF2i3L5,cF2i3L5,F2i3L5_inp1,F2i3L5_inp2,F2i3L5_inp3 );

wire F1i3L6_inp1, F1i3L6_inp2, F1i3L6_inp3;
assign F1i3L6_inp1 = PP[5][1];
assign F1i3L6_inp2 = PP[6][0];
assign F1i3L6_inp3 = C[6];
wire sF1i3L6, cF1i3L6;
FA F1i3L6( sF1i3L6,cF1i3L6,F1i3L6_inp1,F1i3L6_inp2,F1i3L6_inp3 );

wire F2i3L6_inp1, F2i3L6_inp2, F2i3L6_inp3;
assign F2i3L6_inp1 = cHi2L5;
assign F2i3L6_inp2 = sF1i2L6;
assign F2i3L6_inp3 = sHi2L6;
wire sF2i3L6, cF2i3L6;
FA F2i3L6( sF2i3L6,cF2i3L6,F2i3L6_inp1,F2i3L6_inp2,F2i3L6_inp3 );

wire F1i3L7_inp1, F1i3L7_inp2, F1i3L7_inp3;
assign F1i3L7_inp1 = C[7];
assign F1i3L7_inp2 = cF1i2L6;
assign F1i3L7_inp3 = cHi2L6;
wire sF1i3L7, cF1i3L7;
FA F1i3L7( sF1i3L7,cF1i3L7,F1i3L7_inp1,F1i3L7_inp2,F1i3L7_inp3 );

wire F2i3L7_inp1, F2i3L7_inp2, F2i3L7_inp3;
assign F2i3L7_inp1 = sF1i2L7;
assign F2i3L7_inp2 = sF2i2L7;
assign F2i3L7_inp3 = sHi2L7;
wire sF2i3L7, cF2i3L7;
FA F2i3L7( sF2i3L7,cF2i3L7,F2i3L7_inp1,F2i3L7_inp2,F2i3L7_inp3 );

wire F1i3L8_inp1, F1i3L8_inp2, F1i3L8_inp3;
assign F1i3L8_inp1 = cF1i2L7;
assign F1i3L8_inp2 = cF2i2L7;
assign F1i3L8_inp3 = cHi2L7;
wire sF1i3L8, cF1i3L8;
FA F1i3L8( sF1i3L8,cF1i3L8,F1i3L8_inp1,F1i3L8_inp2,F1i3L8_inp3 );

wire F2i3L8_inp1, F2i3L8_inp2, F2i3L8_inp3;
assign F2i3L8_inp1 = sF1i2L8;
assign F2i3L8_inp2 = sF2i2L8;
assign F2i3L8_inp3 = sF3i2L8;
wire sF2i3L8, cF2i3L8;
FA F2i3L8( sF2i3L8,cF2i3L8,F2i3L8_inp1,F2i3L8_inp2,F2i3L8_inp3 );

wire F1i3L9_inp1, F1i3L9_inp2, F1i3L9_inp3;
assign F1i3L9_inp1 = cF1i2L8;
assign F1i3L9_inp2 = cF2i2L8;
assign F1i3L9_inp3 = cF3i2L8;
wire sF1i3L9, cF1i3L9;
FA F1i3L9( sF1i3L9,cF1i3L9,F1i3L9_inp1,F1i3L9_inp2,F1i3L9_inp3 );

wire F2i3L9_inp1, F2i3L9_inp2, F2i3L9_inp3;
assign F2i3L9_inp1 = sF1i2L9;
assign F2i3L9_inp2 = sF2i2L9;
assign F2i3L9_inp3 = sF3i2L9;
wire sF2i3L9, cF2i3L9;
FA F2i3L9( sF2i3L9,cF2i3L9,F2i3L9_inp1,F2i3L9_inp2,F2i3L9_inp3 );

wire F1i3L10_inp1, F1i3L10_inp2, F1i3L10_inp3;
assign F1i3L10_inp1 = cF1i2L9;
assign F1i3L10_inp2 = cF2i2L9;
assign F1i3L10_inp3 = cF3i2L9;
wire sF1i3L10, cF1i3L10;
FA F1i3L10( sF1i3L10,cF1i3L10,F1i3L10_inp1,F1i3L10_inp2,F1i3L10_inp3 );

wire F2i3L10_inp1, F2i3L10_inp2, F2i3L10_inp3;
assign F2i3L10_inp1 = sF1i2L10;
assign F2i3L10_inp2 = sF2i2L10;
assign F2i3L10_inp3 = sF3i2L10;
wire sF2i3L10, cF2i3L10;
FA F2i3L10( sF2i3L10,cF2i3L10,F2i3L10_inp1,F2i3L10_inp2,F2i3L10_inp3 );

wire F1i3L11_inp1, F1i3L11_inp2, F1i3L11_inp3;
assign F1i3L11_inp1 = cF1i2L10;
assign F1i3L11_inp2 = cF2i2L10;
assign F1i3L11_inp3 = cF3i2L10;
wire sF1i3L11, cF1i3L11;
FA F1i3L11( sF1i3L11,cF1i3L11,F1i3L11_inp1,F1i3L11_inp2,F1i3L11_inp3 );

wire F2i3L11_inp1, F2i3L11_inp2, F2i3L11_inp3;
assign F2i3L11_inp1 = sF1i2L11;
assign F2i3L11_inp2 = sF2i2L11;
assign F2i3L11_inp3 = sF3i2L11;
wire sF2i3L11, cF2i3L11;
FA F2i3L11( sF2i3L11,cF2i3L11,F2i3L11_inp1,F2i3L11_inp2,F2i3L11_inp3 );

wire F1i3L12_inp1, F1i3L12_inp2, F1i3L12_inp3;
assign F1i3L12_inp1 = cF1i2L11;
assign F1i3L12_inp2 = cF2i2L11;
assign F1i3L12_inp3 = cF3i2L11;
wire sF1i3L12, cF1i3L12;
FA F1i3L12( sF1i3L12,cF1i3L12,F1i3L12_inp1,F1i3L12_inp2,F1i3L12_inp3 );

wire F2i3L12_inp1, F2i3L12_inp2, F2i3L12_inp3;
assign F2i3L12_inp1 = sF1i2L12;
assign F2i3L12_inp2 = sF2i2L12;
assign F2i3L12_inp3 = sF3i2L12;
wire sF2i3L12, cF2i3L12;
FA F2i3L12( sF2i3L12,cF2i3L12,F2i3L12_inp1,F2i3L12_inp2,F2i3L12_inp3 );

wire F1i3L13_inp1, F1i3L13_inp2, F1i3L13_inp3;
assign F1i3L13_inp1 = cF1i2L12;
assign F1i3L13_inp2 = cF2i2L12;
assign F1i3L13_inp3 = cF3i2L12;
wire sF1i3L13, cF1i3L13;
FA F1i3L13( sF1i3L13,cF1i3L13,F1i3L13_inp1,F1i3L13_inp2,F1i3L13_inp3 );

wire F2i3L13_inp1, F2i3L13_inp2, F2i3L13_inp3;
assign F2i3L13_inp1 = sF1i2L13;
assign F2i3L13_inp2 = sF2i2L13;
assign F2i3L13_inp3 = sF3i2L13;
wire sF2i3L13, cF2i3L13;
FA F2i3L13( sF2i3L13,cF2i3L13,F2i3L13_inp1,F2i3L13_inp2,F2i3L13_inp3 );

wire F1i3L14_inp1, F1i3L14_inp2, F1i3L14_inp3;
assign F1i3L14_inp1 = PP[10][4];
assign F1i3L14_inp2 = cF1i2L13;
assign F1i3L14_inp3 = cF2i2L13;
wire sF1i3L14, cF1i3L14;
FA F1i3L14( sF1i3L14,cF1i3L14,F1i3L14_inp1,F1i3L14_inp2,F1i3L14_inp3 );

wire F2i3L14_inp1, F2i3L14_inp2, F2i3L14_inp3;
assign F2i3L14_inp1 = cF3i2L13;
assign F2i3L14_inp2 = sF1i2L14;
assign F2i3L14_inp3 = sF2i2L14;
wire sF2i3L14, cF2i3L14;
FA F2i3L14( sF2i3L14,cF2i3L14,F2i3L14_inp1,F2i3L14_inp2,F2i3L14_inp3 );

wire F1i3L15_inp1, F1i3L15_inp2, F1i3L15_inp3;
assign F1i3L15_inp1 = PP[8][7];
assign F1i3L15_inp2 = PP[9][6];
assign F1i3L15_inp3 = PP[10][5];
wire sF1i3L15, cF1i3L15;
FA F1i3L15( sF1i3L15,cF1i3L15,F1i3L15_inp1,F1i3L15_inp2,F1i3L15_inp3 );

wire F2i3L15_inp1, F2i3L15_inp2, F2i3L15_inp3;
assign F2i3L15_inp1 = cF1i2L14;
assign F2i3L15_inp2 = cF2i2L14;
assign F2i3L15_inp3 = sF1i2L15;
wire sF2i3L15, cF2i3L15;
FA F2i3L15( sF2i3L15,cF2i3L15,F2i3L15_inp1,F2i3L15_inp2,F2i3L15_inp3 );

wire F1i3L16_inp1, F1i3L16_inp2, F1i3L16_inp3;
assign F1i3L16_inp1 = PP[6][10];
assign F1i3L16_inp2 = PP[7][9];
assign F1i3L16_inp3 = PP[8][8];
wire sF1i3L16, cF1i3L16;
FA F1i3L16( sF1i3L16,cF1i3L16,F1i3L16_inp1,F1i3L16_inp2,F1i3L16_inp3 );

wire F2i3L16_inp1, F2i3L16_inp2, F2i3L16_inp3;
assign F2i3L16_inp1 = PP[9][7];
assign F2i3L16_inp2 = PP[10][6];
assign F2i3L16_inp3 = cF1i2L15;
wire sF2i3L16, cF2i3L16;
FA F2i3L16( sF2i3L16,cF2i3L16,F2i3L16_inp1,F2i3L16_inp2,F2i3L16_inp3 );

wire F1i3L17_inp1, F1i3L17_inp2, F1i3L17_inp3;
assign F1i3L17_inp1 = PP[7][10];
assign F1i3L17_inp2 = PP[8][9];
assign F1i3L17_inp3 = PP[9][8];
wire sF1i3L17, cF1i3L17;
FA F1i3L17( sF1i3L17,cF1i3L17,F1i3L17_inp1,F1i3L17_inp2,F1i3L17_inp3 );



///////////// Iteration Number =4///////////////////





wire Hi4L2_inp1, Hi4L2_inp2;
assign Hi4L2_inp1 = PP[0][2];
assign Hi4L2_inp2 = PP[1][1];
wire sHi4L2, cHi4L2;
HA Hi4L2 ( sHi4L2,cHi4L2,Hi4L2_inp1,Hi4L2_inp2 );

wire F1i4L3_inp1, F1i4L3_inp2, F1i4L3_inp3;
assign F1i4L3_inp1 = PP[2][1];
assign F1i4L3_inp2 = PP[3][0];
assign F1i4L3_inp3 = C[3];
wire sF1i4L3, cF1i4L3;
FA F1i4L3( sF1i4L3,cF1i4L3,F1i4L3_inp1,F1i4L3_inp2,F1i4L3_inp3 );

wire F1i4L4_inp1, F1i4L4_inp2, F1i4L4_inp3;
assign F1i4L4_inp1 = C[4];
assign F1i4L4_inp2 = cHi3L3;
assign F1i4L4_inp3 = sF1i3L4;
wire sF1i4L4, cF1i4L4;
FA F1i4L4( sF1i4L4,cF1i4L4,F1i4L4_inp1,F1i4L4_inp2,F1i4L4_inp3 );

wire F1i4L5_inp1, F1i4L5_inp2, F1i4L5_inp3;
assign F1i4L5_inp1 = cF1i3L4;
assign F1i4L5_inp2 = cHi3L4;
assign F1i4L5_inp3 = sF1i3L5;
wire sF1i4L5, cF1i4L5;
FA F1i4L5( sF1i4L5,cF1i4L5,F1i4L5_inp1,F1i4L5_inp2,F1i4L5_inp3 );

wire F1i4L6_inp1, F1i4L6_inp2, F1i4L6_inp3;
assign F1i4L6_inp1 = cF1i3L5;
assign F1i4L6_inp2 = cF2i3L5;
assign F1i4L6_inp3 = sF1i3L6;
wire sF1i4L6, cF1i4L6;
FA F1i4L6( sF1i4L6,cF1i4L6,F1i4L6_inp1,F1i4L6_inp2,F1i4L6_inp3 );

wire F1i4L7_inp1, F1i4L7_inp2, F1i4L7_inp3;
assign F1i4L7_inp1 = cF1i3L6;
assign F1i4L7_inp2 = cF2i3L6;
assign F1i4L7_inp3 = sF1i3L7;
wire sF1i4L7, cF1i4L7;
FA F1i4L7( sF1i4L7,cF1i4L7,F1i4L7_inp1,F1i4L7_inp2,F1i4L7_inp3 );

wire F1i4L8_inp1, F1i4L8_inp2, F1i4L8_inp3;
assign F1i4L8_inp1 = cF1i3L7;
assign F1i4L8_inp2 = cF2i3L7;
assign F1i4L8_inp3 = sF1i3L8;
wire sF1i4L8, cF1i4L8;
FA F1i4L8( sF1i4L8,cF1i4L8,F1i4L8_inp1,F1i4L8_inp2,F1i4L8_inp3 );

wire F1i4L9_inp1, F1i4L9_inp2, F1i4L9_inp3;
assign F1i4L9_inp1 = cF1i3L8;
assign F1i4L9_inp2 = cF2i3L8;
assign F1i4L9_inp3 = sF1i3L9;
wire sF1i4L9, cF1i4L9;
FA F1i4L9( sF1i4L9,cF1i4L9,F1i4L9_inp1,F1i4L9_inp2,F1i4L9_inp3 );

wire F1i4L10_inp1, F1i4L10_inp2, F1i4L10_inp3;
assign F1i4L10_inp1 = cF1i3L9;
assign F1i4L10_inp2 = cF2i3L9;
assign F1i4L10_inp3 = sF1i3L10;
wire sF1i4L10, cF1i4L10;
FA F1i4L10( sF1i4L10,cF1i4L10,F1i4L10_inp1,F1i4L10_inp2,F1i4L10_inp3 );

wire F1i4L11_inp1, F1i4L11_inp2, F1i4L11_inp3;
assign F1i4L11_inp1 = cF1i3L10;
assign F1i4L11_inp2 = cF2i3L10;
assign F1i4L11_inp3 = sF1i3L11;
wire sF1i4L11, cF1i4L11;
FA F1i4L11( sF1i4L11,cF1i4L11,F1i4L11_inp1,F1i4L11_inp2,F1i4L11_inp3 );

wire F1i4L12_inp1, F1i4L12_inp2, F1i4L12_inp3;
assign F1i4L12_inp1 = cF1i3L11;
assign F1i4L12_inp2 = cF2i3L11;
assign F1i4L12_inp3 = sF1i3L12;
wire sF1i4L12, cF1i4L12;
FA F1i4L12( sF1i4L12,cF1i4L12,F1i4L12_inp1,F1i4L12_inp2,F1i4L12_inp3 );

wire F1i4L13_inp1, F1i4L13_inp2, F1i4L13_inp3;
assign F1i4L13_inp1 = cF1i3L12;
assign F1i4L13_inp2 = cF2i3L12;
assign F1i4L13_inp3 = sF1i3L13;
wire sF1i4L13, cF1i4L13;
FA F1i4L13( sF1i4L13,cF1i4L13,F1i4L13_inp1,F1i4L13_inp2,F1i4L13_inp3 );

wire F1i4L14_inp1, F1i4L14_inp2, F1i4L14_inp3;
assign F1i4L14_inp1 = cF1i3L13;
assign F1i4L14_inp2 = cF2i3L13;
assign F1i4L14_inp3 = sF1i3L14;
wire sF1i4L14, cF1i4L14;
FA F1i4L14( sF1i4L14,cF1i4L14,F1i4L14_inp1,F1i4L14_inp2,F1i4L14_inp3 );

wire F1i4L15_inp1, F1i4L15_inp2, F1i4L15_inp3;
assign F1i4L15_inp1 = cF1i3L14;
assign F1i4L15_inp2 = cF2i3L14;
assign F1i4L15_inp3 = sF1i3L15;
wire sF1i4L15, cF1i4L15;
FA F1i4L15( sF1i4L15,cF1i4L15,F1i4L15_inp1,F1i4L15_inp2,F1i4L15_inp3 );

wire F1i4L16_inp1, F1i4L16_inp2, F1i4L16_inp3;
assign F1i4L16_inp1 = cF1i3L15;
assign F1i4L16_inp2 = cF2i3L15;
assign F1i4L16_inp3 = sF1i3L16;
wire sF1i4L16, cF1i4L16;
FA F1i4L16( sF1i4L16,cF1i4L16,F1i4L16_inp1,F1i4L16_inp2,F1i4L16_inp3 );

wire F1i4L17_inp1, F1i4L17_inp2, F1i4L17_inp3;
assign F1i4L17_inp1 = PP[10][7];
assign F1i4L17_inp2 = cF1i3L16;
assign F1i4L17_inp3 = cF2i3L16;
wire sF1i4L17, cF1i4L17;
FA F1i4L17( sF1i4L17,cF1i4L17,F1i4L17_inp1,F1i4L17_inp2,F1i4L17_inp3 );

wire F1i4L18_inp1, F1i4L18_inp2, F1i4L18_inp3;
assign F1i4L18_inp1 = PP[8][10];
assign F1i4L18_inp2 = PP[9][9];
assign F1i4L18_inp3 = PP[10][8];
wire sF1i4L18, cF1i4L18;
FA F1i4L18( sF1i4L18,cF1i4L18,F1i4L18_inp1,F1i4L18_inp2,F1i4L18_inp3 );



///////////// Iteration Number =5///////////////////





wire Hi5L1_inp1, Hi5L1_inp2;
assign Hi5L1_inp1 = PP[0][1];
assign Hi5L1_inp2 = PP[1][0];
wire sHi5L1, cHi5L1;
HA Hi5L1 ( sHi5L1,cHi5L1,Hi5L1_inp1,Hi5L1_inp2 );

wire F1i5L2_inp1, F1i5L2_inp2, F1i5L2_inp3;
assign F1i5L2_inp1 = PP[2][0];
assign F1i5L2_inp2 = C[2];
assign F1i5L2_inp3 = sHi4L2;
wire sF1i5L2, cF1i5L2;
FA F1i5L2( sF1i5L2,cF1i5L2,F1i5L2_inp1,F1i5L2_inp2,F1i5L2_inp3 );

wire F1i5L3_inp1, F1i5L3_inp2, F1i5L3_inp3;
assign F1i5L3_inp1 = sHi3L3;
assign F1i5L3_inp2 = cHi4L2;
assign F1i5L3_inp3 = sF1i4L3;
wire sF1i5L3, cF1i5L3;
FA F1i5L3( sF1i5L3,cF1i5L3,F1i5L3_inp1,F1i5L3_inp2,F1i5L3_inp3 );

wire F1i5L4_inp1, F1i5L4_inp2, F1i5L4_inp3;
assign F1i5L4_inp1 = sHi3L4;
assign F1i5L4_inp2 = cF1i4L3;
assign F1i5L4_inp3 = sF1i4L4;
wire sF1i5L4, cF1i5L4;
FA F1i5L4( sF1i5L4,cF1i5L4,F1i5L4_inp1,F1i5L4_inp2,F1i5L4_inp3 );

wire F1i5L5_inp1, F1i5L5_inp2, F1i5L5_inp3;
assign F1i5L5_inp1 = sF2i3L5;
assign F1i5L5_inp2 = cF1i4L4;
assign F1i5L5_inp3 = sF1i4L5;
wire sF1i5L5, cF1i5L5;
FA F1i5L5( sF1i5L5,cF1i5L5,F1i5L5_inp1,F1i5L5_inp2,F1i5L5_inp3 );

wire F1i5L6_inp1, F1i5L6_inp2, F1i5L6_inp3;
assign F1i5L6_inp1 = sF2i3L6;
assign F1i5L6_inp2 = cF1i4L5;
assign F1i5L6_inp3 = sF1i4L6;
wire sF1i5L6, cF1i5L6;
FA F1i5L6( sF1i5L6,cF1i5L6,F1i5L6_inp1,F1i5L6_inp2,F1i5L6_inp3 );

wire F1i5L7_inp1, F1i5L7_inp2, F1i5L7_inp3;
assign F1i5L7_inp1 = sF2i3L7;
assign F1i5L7_inp2 = cF1i4L6;
assign F1i5L7_inp3 = sF1i4L7;
wire sF1i5L7, cF1i5L7;
FA F1i5L7( sF1i5L7,cF1i5L7,F1i5L7_inp1,F1i5L7_inp2,F1i5L7_inp3 );

wire F1i5L8_inp1, F1i5L8_inp2, F1i5L8_inp3;
assign F1i5L8_inp1 = sF2i3L8;
assign F1i5L8_inp2 = cF1i4L7;
assign F1i5L8_inp3 = sF1i4L8;
wire sF1i5L8, cF1i5L8;
FA F1i5L8( sF1i5L8,cF1i5L8,F1i5L8_inp1,F1i5L8_inp2,F1i5L8_inp3 );

wire F1i5L9_inp1, F1i5L9_inp2, F1i5L9_inp3;
assign F1i5L9_inp1 = sF2i3L9;
assign F1i5L9_inp2 = cF1i4L8;
assign F1i5L9_inp3 = sF1i4L9;
wire sF1i5L9, cF1i5L9;
FA F1i5L9( sF1i5L9,cF1i5L9,F1i5L9_inp1,F1i5L9_inp2,F1i5L9_inp3 );

wire F1i5L10_inp1, F1i5L10_inp2, F1i5L10_inp3;
assign F1i5L10_inp1 = sF2i3L10;
assign F1i5L10_inp2 = cF1i4L9;
assign F1i5L10_inp3 = sF1i4L10;
wire sF1i5L10, cF1i5L10;
FA F1i5L10( sF1i5L10,cF1i5L10,F1i5L10_inp1,F1i5L10_inp2,F1i5L10_inp3 );

wire F1i5L11_inp1, F1i5L11_inp2, F1i5L11_inp3;
assign F1i5L11_inp1 = sF2i3L11;
assign F1i5L11_inp2 = cF1i4L10;
assign F1i5L11_inp3 = sF1i4L11;
wire sF1i5L11, cF1i5L11;
FA F1i5L11( sF1i5L11,cF1i5L11,F1i5L11_inp1,F1i5L11_inp2,F1i5L11_inp3 );

wire F1i5L12_inp1, F1i5L12_inp2, F1i5L12_inp3;
assign F1i5L12_inp1 = sF2i3L12;
assign F1i5L12_inp2 = cF1i4L11;
assign F1i5L12_inp3 = sF1i4L12;
wire sF1i5L12, cF1i5L12;
FA F1i5L12( sF1i5L12,cF1i5L12,F1i5L12_inp1,F1i5L12_inp2,F1i5L12_inp3 );

wire F1i5L13_inp1, F1i5L13_inp2, F1i5L13_inp3;
assign F1i5L13_inp1 = sF2i3L13;
assign F1i5L13_inp2 = cF1i4L12;
assign F1i5L13_inp3 = sF1i4L13;
wire sF1i5L13, cF1i5L13;
FA F1i5L13( sF1i5L13,cF1i5L13,F1i5L13_inp1,F1i5L13_inp2,F1i5L13_inp3 );

wire F1i5L14_inp1, F1i5L14_inp2, F1i5L14_inp3;
assign F1i5L14_inp1 = sF2i3L14;
assign F1i5L14_inp2 = cF1i4L13;
assign F1i5L14_inp3 = sF1i4L14;
wire sF1i5L14, cF1i5L14;
FA F1i5L14( sF1i5L14,cF1i5L14,F1i5L14_inp1,F1i5L14_inp2,F1i5L14_inp3 );

wire F1i5L15_inp1, F1i5L15_inp2, F1i5L15_inp3;
assign F1i5L15_inp1 = sF2i3L15;
assign F1i5L15_inp2 = cF1i4L14;
assign F1i5L15_inp3 = sF1i4L15;
wire sF1i5L15, cF1i5L15;
FA F1i5L15( sF1i5L15,cF1i5L15,F1i5L15_inp1,F1i5L15_inp2,F1i5L15_inp3 );

wire F1i5L16_inp1, F1i5L16_inp2, F1i5L16_inp3;
assign F1i5L16_inp1 = sF2i3L16;
assign F1i5L16_inp2 = cF1i4L15;
assign F1i5L16_inp3 = sF1i4L16;
wire sF1i5L16, cF1i5L16;
FA F1i5L16( sF1i5L16,cF1i5L16,F1i5L16_inp1,F1i5L16_inp2,F1i5L16_inp3 );

wire F1i5L17_inp1, F1i5L17_inp2, F1i5L17_inp3;
assign F1i5L17_inp1 = sF1i3L17;
assign F1i5L17_inp2 = cF1i4L16;
assign F1i5L17_inp3 = sF1i4L17;
wire sF1i5L17, cF1i5L17;
FA F1i5L17( sF1i5L17,cF1i5L17,F1i5L17_inp1,F1i5L17_inp2,F1i5L17_inp3 );

wire F1i5L18_inp1, F1i5L18_inp2, F1i5L18_inp3;
assign F1i5L18_inp1 = cF1i3L17;
assign F1i5L18_inp2 = cF1i4L17;
assign F1i5L18_inp3 = sF1i4L18;
wire sF1i5L18, cF1i5L18;
FA F1i5L18( sF1i5L18,cF1i5L18,F1i5L18_inp1,F1i5L18_inp2,F1i5L18_inp3 );

wire F1i5L19_inp1, F1i5L19_inp2, F1i5L19_inp3;
assign F1i5L19_inp1 = PP[9][10];
assign F1i5L19_inp2 = PP[10][9];
assign F1i5L19_inp3 = cF1i4L18;
wire sF1i5L19, cF1i5L19;
FA F1i5L19( sF1i5L19,cF1i5L19,F1i5L19_inp1,F1i5L19_inp2,F1i5L19_inp3 );


assign out1 ={{1'b0},{PP[10][10]},{cF1i5L18},{cF1i5L17},{cF1i5L16},{cF1i5L15},{cF1i5L14},{cF1i5L13},{cF1i5L12},{cF1i5L11},{cF1i5L10},{cF1i5L9},{cF1i5L8},{cF1i5L7},{cF1i5L6},{cF1i5L5},{cF1i5L4},{cF1i5L3},{cF1i5L2},{cHi5L1},{C[1]},{PP[0][0]}};
assign out2 ={{1'b0},{cF1i5L19},{sF1i5L19},{sF1i5L18},{sF1i5L17},{sF1i5L16},{sF1i5L15},{sF1i5L14},{sF1i5L13},{sF1i5L12},{sF1i5L11},{sF1i5L10},{sF1i5L9},{sF1i5L8},{sF1i5L7},{sF1i5L6},{sF1i5L5},{sF1i5L4},{sF1i5L3},{sF1i5L2},{sHi5L1},{C[0]}} ;
endmodule