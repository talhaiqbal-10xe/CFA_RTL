module adder8x12(
output [14:0] out1,out2,
input [11:0]A,B,C,D,E,F,G,H );


wire [14:0] CV;
 assign CV=15'b000000000000100;




///////////// Iteration Number =1///////////////////





wire F1i1L0_inp1, F1i1L0_inp2, F1i1L0_inp3;
assign F1i1L0_inp1 = A[0];
assign F1i1L0_inp2 = B[0];
assign F1i1L0_inp3 = C[0];
wire sF1i1L0, cF1i1L0;
FA F1i1L0( sF1i1L0,cF1i1L0,F1i1L0_inp1,F1i1L0_inp2,F1i1L0_inp3 );

wire F1i1L1_inp1, F1i1L1_inp2, F1i1L1_inp3;
assign F1i1L1_inp1 = A[1];
assign F1i1L1_inp2 = B[1];
assign F1i1L1_inp3 = C[1];
wire sF1i1L1, cF1i1L1;
FA F1i1L1( sF1i1L1,cF1i1L1,F1i1L1_inp1,F1i1L1_inp2,F1i1L1_inp3 );

wire Hi1L1_inp1, Hi1L1_inp2;
assign Hi1L1_inp1 = D[1];
assign Hi1L1_inp2 = E[1];
wire sHi1L1, cHi1L1;
HA Hi1L1 ( sHi1L1,cHi1L1,Hi1L1_inp1,Hi1L1_inp2 );

wire F1i1L2_inp1, F1i1L2_inp2, F1i1L2_inp3;
assign F1i1L2_inp1 = A[2];
assign F1i1L2_inp2 = B[2];
assign F1i1L2_inp3 = C[2];
wire sF1i1L2, cF1i1L2;
FA F1i1L2( sF1i1L2,cF1i1L2,F1i1L2_inp1,F1i1L2_inp2,F1i1L2_inp3 );

wire F2i1L2_inp1, F2i1L2_inp2, F2i1L2_inp3;
assign F2i1L2_inp1 = D[2];
assign F2i1L2_inp2 = E[2];
assign F2i1L2_inp3 = F[2];
wire sF2i1L2, cF2i1L2;
FA F2i1L2( sF2i1L2,cF2i1L2,F2i1L2_inp1,F2i1L2_inp2,F2i1L2_inp3 );

wire Hi1L2_inp1, Hi1L2_inp2;
assign Hi1L2_inp1 = G[2];
assign Hi1L2_inp2 = H[2];
wire sHi1L2, cHi1L2;
HA Hi1L2 ( sHi1L2,cHi1L2,Hi1L2_inp1,Hi1L2_inp2 );

wire F1i1L3_inp1, F1i1L3_inp2, F1i1L3_inp3;
assign F1i1L3_inp1 = A[3];
assign F1i1L3_inp2 = B[3];
assign F1i1L3_inp3 = C[3];
wire sF1i1L3, cF1i1L3;
FA F1i1L3( sF1i1L3,cF1i1L3,F1i1L3_inp1,F1i1L3_inp2,F1i1L3_inp3 );

wire F2i1L3_inp1, F2i1L3_inp2, F2i1L3_inp3;
assign F2i1L3_inp1 = D[3];
assign F2i1L3_inp2 = E[3];
assign F2i1L3_inp3 = F[3];
wire sF2i1L3, cF2i1L3;
FA F2i1L3( sF2i1L3,cF2i1L3,F2i1L3_inp1,F2i1L3_inp2,F2i1L3_inp3 );

wire Hi1L3_inp1, Hi1L3_inp2;
assign Hi1L3_inp1 = G[3];
assign Hi1L3_inp2 = H[3];
wire sHi1L3, cHi1L3;
HA Hi1L3 ( sHi1L3,cHi1L3,Hi1L3_inp1,Hi1L3_inp2 );

wire F1i1L4_inp1, F1i1L4_inp2, F1i1L4_inp3;
assign F1i1L4_inp1 = A[4];
assign F1i1L4_inp2 = B[4];
assign F1i1L4_inp3 = C[4];
wire sF1i1L4, cF1i1L4;
FA F1i1L4( sF1i1L4,cF1i1L4,F1i1L4_inp1,F1i1L4_inp2,F1i1L4_inp3 );

wire F2i1L4_inp1, F2i1L4_inp2, F2i1L4_inp3;
assign F2i1L4_inp1 = D[4];
assign F2i1L4_inp2 = E[4];
assign F2i1L4_inp3 = F[4];
wire sF2i1L4, cF2i1L4;
FA F2i1L4( sF2i1L4,cF2i1L4,F2i1L4_inp1,F2i1L4_inp2,F2i1L4_inp3 );

wire Hi1L4_inp1, Hi1L4_inp2;
assign Hi1L4_inp1 = G[4];
assign Hi1L4_inp2 = H[4];
wire sHi1L4, cHi1L4;
HA Hi1L4 ( sHi1L4,cHi1L4,Hi1L4_inp1,Hi1L4_inp2 );

wire F1i1L5_inp1, F1i1L5_inp2, F1i1L5_inp3;
assign F1i1L5_inp1 = A[5];
assign F1i1L5_inp2 = B[5];
assign F1i1L5_inp3 = C[5];
wire sF1i1L5, cF1i1L5;
FA F1i1L5( sF1i1L5,cF1i1L5,F1i1L5_inp1,F1i1L5_inp2,F1i1L5_inp3 );

wire F2i1L5_inp1, F2i1L5_inp2, F2i1L5_inp3;
assign F2i1L5_inp1 = D[5];
assign F2i1L5_inp2 = E[5];
assign F2i1L5_inp3 = F[5];
wire sF2i1L5, cF2i1L5;
FA F2i1L5( sF2i1L5,cF2i1L5,F2i1L5_inp1,F2i1L5_inp2,F2i1L5_inp3 );

wire Hi1L5_inp1, Hi1L5_inp2;
assign Hi1L5_inp1 = G[5];
assign Hi1L5_inp2 = H[5];
wire sHi1L5, cHi1L5;
HA Hi1L5 ( sHi1L5,cHi1L5,Hi1L5_inp1,Hi1L5_inp2 );

wire F1i1L6_inp1, F1i1L6_inp2, F1i1L6_inp3;
assign F1i1L6_inp1 = A[6];
assign F1i1L6_inp2 = B[6];
assign F1i1L6_inp3 = C[6];
wire sF1i1L6, cF1i1L6;
FA F1i1L6( sF1i1L6,cF1i1L6,F1i1L6_inp1,F1i1L6_inp2,F1i1L6_inp3 );

wire F2i1L6_inp1, F2i1L6_inp2, F2i1L6_inp3;
assign F2i1L6_inp1 = D[6];
assign F2i1L6_inp2 = E[6];
assign F2i1L6_inp3 = F[6];
wire sF2i1L6, cF2i1L6;
FA F2i1L6( sF2i1L6,cF2i1L6,F2i1L6_inp1,F2i1L6_inp2,F2i1L6_inp3 );

wire Hi1L6_inp1, Hi1L6_inp2;
assign Hi1L6_inp1 = G[6];
assign Hi1L6_inp2 = H[6];
wire sHi1L6, cHi1L6;
HA Hi1L6 ( sHi1L6,cHi1L6,Hi1L6_inp1,Hi1L6_inp2 );

wire F1i1L7_inp1, F1i1L7_inp2, F1i1L7_inp3;
assign F1i1L7_inp1 = A[7];
assign F1i1L7_inp2 = B[7];
assign F1i1L7_inp3 = C[7];
wire sF1i1L7, cF1i1L7;
FA F1i1L7( sF1i1L7,cF1i1L7,F1i1L7_inp1,F1i1L7_inp2,F1i1L7_inp3 );

wire F2i1L7_inp1, F2i1L7_inp2, F2i1L7_inp3;
assign F2i1L7_inp1 = D[7];
assign F2i1L7_inp2 = E[7];
assign F2i1L7_inp3 = F[7];
wire sF2i1L7, cF2i1L7;
FA F2i1L7( sF2i1L7,cF2i1L7,F2i1L7_inp1,F2i1L7_inp2,F2i1L7_inp3 );

wire Hi1L7_inp1, Hi1L7_inp2;
assign Hi1L7_inp1 = G[7];
assign Hi1L7_inp2 = H[7];
wire sHi1L7, cHi1L7;
HA Hi1L7 ( sHi1L7,cHi1L7,Hi1L7_inp1,Hi1L7_inp2 );

wire F1i1L8_inp1, F1i1L8_inp2, F1i1L8_inp3;
assign F1i1L8_inp1 = A[8];
assign F1i1L8_inp2 = B[8];
assign F1i1L8_inp3 = C[8];
wire sF1i1L8, cF1i1L8;
FA F1i1L8( sF1i1L8,cF1i1L8,F1i1L8_inp1,F1i1L8_inp2,F1i1L8_inp3 );

wire F2i1L8_inp1, F2i1L8_inp2, F2i1L8_inp3;
assign F2i1L8_inp1 = D[8];
assign F2i1L8_inp2 = E[8];
assign F2i1L8_inp3 = F[8];
wire sF2i1L8, cF2i1L8;
FA F2i1L8( sF2i1L8,cF2i1L8,F2i1L8_inp1,F2i1L8_inp2,F2i1L8_inp3 );

wire Hi1L8_inp1, Hi1L8_inp2;
assign Hi1L8_inp1 = G[8];
assign Hi1L8_inp2 = H[8];
wire sHi1L8, cHi1L8;
HA Hi1L8 ( sHi1L8,cHi1L8,Hi1L8_inp1,Hi1L8_inp2 );

wire F1i1L9_inp1, F1i1L9_inp2, F1i1L9_inp3;
assign F1i1L9_inp1 = A[9];
assign F1i1L9_inp2 = B[9];
assign F1i1L9_inp3 = C[9];
wire sF1i1L9, cF1i1L9;
FA F1i1L9( sF1i1L9,cF1i1L9,F1i1L9_inp1,F1i1L9_inp2,F1i1L9_inp3 );

wire F2i1L9_inp1, F2i1L9_inp2, F2i1L9_inp3;
assign F2i1L9_inp1 = D[9];
assign F2i1L9_inp2 = E[9];
assign F2i1L9_inp3 = F[9];
wire sF2i1L9, cF2i1L9;
FA F2i1L9( sF2i1L9,cF2i1L9,F2i1L9_inp1,F2i1L9_inp2,F2i1L9_inp3 );

wire Hi1L9_inp1, Hi1L9_inp2;
assign Hi1L9_inp1 = G[9];
assign Hi1L9_inp2 = H[9];
wire sHi1L9, cHi1L9;
HA Hi1L9 ( sHi1L9,cHi1L9,Hi1L9_inp1,Hi1L9_inp2 );

wire F1i1L10_inp1, F1i1L10_inp2, F1i1L10_inp3;
assign F1i1L10_inp1 = A[10];
assign F1i1L10_inp2 = B[10];
assign F1i1L10_inp3 = C[10];
wire sF1i1L10, cF1i1L10;
FA F1i1L10( sF1i1L10,cF1i1L10,F1i1L10_inp1,F1i1L10_inp2,F1i1L10_inp3 );

wire F2i1L10_inp1, F2i1L10_inp2, F2i1L10_inp3;
assign F2i1L10_inp1 = D[10];
assign F2i1L10_inp2 = E[10];
assign F2i1L10_inp3 = F[10];
wire sF2i1L10, cF2i1L10;
FA F2i1L10( sF2i1L10,cF2i1L10,F2i1L10_inp1,F2i1L10_inp2,F2i1L10_inp3 );

wire Hi1L10_inp1, Hi1L10_inp2;
assign Hi1L10_inp1 = G[10];
assign Hi1L10_inp2 = H[10];
wire sHi1L10, cHi1L10;
HA Hi1L10 ( sHi1L10,cHi1L10,Hi1L10_inp1,Hi1L10_inp2 );

wire F1i1L11_inp1, F1i1L11_inp2, F1i1L11_inp3;
assign F1i1L11_inp1 = A[11];
assign F1i1L11_inp2 = B[11];
assign F1i1L11_inp3 = C[11];
wire sF1i1L11, cF1i1L11;
FA F1i1L11( sF1i1L11,cF1i1L11,F1i1L11_inp1,F1i1L11_inp2,F1i1L11_inp3 );

wire F2i1L11_inp1, F2i1L11_inp2, F2i1L11_inp3;
assign F2i1L11_inp1 = D[11];
assign F2i1L11_inp2 = E[11];
assign F2i1L11_inp3 = F[11];
wire sF2i1L11, cF2i1L11;
FA F2i1L11( sF2i1L11,cF2i1L11,F2i1L11_inp1,F2i1L11_inp2,F2i1L11_inp3 );

wire Hi1L11_inp1, Hi1L11_inp2;
assign Hi1L11_inp1 = G[11];
assign Hi1L11_inp2 = H[11];
wire sHi1L11, cHi1L11;
HA Hi1L11 ( sHi1L11,cHi1L11,Hi1L11_inp1,Hi1L11_inp2 );



///////////// Iteration Number =2///////////////////





wire F1i2L0_inp1, F1i2L0_inp2, F1i2L0_inp3;
assign F1i2L0_inp1 = D[0];
assign F1i2L0_inp2 = E[0];
assign F1i2L0_inp3 = F[0];
wire sF1i2L0, cF1i2L0;
FA F1i2L0( sF1i2L0,cF1i2L0,F1i2L0_inp1,F1i2L0_inp2,F1i2L0_inp3 );

wire F1i2L1_inp1, F1i2L1_inp2, F1i2L1_inp3;
assign F1i2L1_inp1 = F[1];
assign F1i2L1_inp2 = G[1];
assign F1i2L1_inp3 = H[1];
wire sF1i2L1, cF1i2L1;
FA F1i2L1( sF1i2L1,cF1i2L1,F1i2L1_inp1,F1i2L1_inp2,F1i2L1_inp3 );

wire Hi2L1_inp1, Hi2L1_inp2;
assign Hi2L1_inp1 = cF1i1L0;
assign Hi2L1_inp2 = sF1i1L1;
wire sHi2L1, cHi2L1;
HA Hi2L1 ( sHi2L1,cHi2L1,Hi2L1_inp1,Hi2L1_inp2 );

wire F1i2L2_inp1, F1i2L2_inp2, F1i2L2_inp3;
assign F1i2L2_inp1 = CV[2];
assign F1i2L2_inp2 = cF1i1L1;
assign F1i2L2_inp3 = cHi1L1;
wire sF1i2L2, cF1i2L2;
FA F1i2L2( sF1i2L2,cF1i2L2,F1i2L2_inp1,F1i2L2_inp2,F1i2L2_inp3 );

wire F2i2L2_inp1, F2i2L2_inp2, F2i2L2_inp3;
assign F2i2L2_inp1 = sF1i1L2;
assign F2i2L2_inp2 = sF2i1L2;
assign F2i2L2_inp3 = sHi1L2;
wire sF2i2L2, cF2i2L2;
FA F2i2L2( sF2i2L2,cF2i2L2,F2i2L2_inp1,F2i2L2_inp2,F2i2L2_inp3 );

wire F1i2L3_inp1, F1i2L3_inp2, F1i2L3_inp3;
assign F1i2L3_inp1 = cF1i1L2;
assign F1i2L3_inp2 = cF2i1L2;
assign F1i2L3_inp3 = cHi1L2;
wire sF1i2L3, cF1i2L3;
FA F1i2L3( sF1i2L3,cF1i2L3,F1i2L3_inp1,F1i2L3_inp2,F1i2L3_inp3 );

wire F2i2L3_inp1, F2i2L3_inp2, F2i2L3_inp3;
assign F2i2L3_inp1 = sF1i1L3;
assign F2i2L3_inp2 = sF2i1L3;
assign F2i2L3_inp3 = sHi1L3;
wire sF2i2L3, cF2i2L3;
FA F2i2L3( sF2i2L3,cF2i2L3,F2i2L3_inp1,F2i2L3_inp2,F2i2L3_inp3 );

wire F1i2L4_inp1, F1i2L4_inp2, F1i2L4_inp3;
assign F1i2L4_inp1 = cF1i1L3;
assign F1i2L4_inp2 = cF2i1L3;
assign F1i2L4_inp3 = cHi1L3;
wire sF1i2L4, cF1i2L4;
FA F1i2L4( sF1i2L4,cF1i2L4,F1i2L4_inp1,F1i2L4_inp2,F1i2L4_inp3 );

wire F2i2L4_inp1, F2i2L4_inp2, F2i2L4_inp3;
assign F2i2L4_inp1 = sF1i1L4;
assign F2i2L4_inp2 = sF2i1L4;
assign F2i2L4_inp3 = sHi1L4;
wire sF2i2L4, cF2i2L4;
FA F2i2L4( sF2i2L4,cF2i2L4,F2i2L4_inp1,F2i2L4_inp2,F2i2L4_inp3 );

wire F1i2L5_inp1, F1i2L5_inp2, F1i2L5_inp3;
assign F1i2L5_inp1 = cF1i1L4;
assign F1i2L5_inp2 = cF2i1L4;
assign F1i2L5_inp3 = cHi1L4;
wire sF1i2L5, cF1i2L5;
FA F1i2L5( sF1i2L5,cF1i2L5,F1i2L5_inp1,F1i2L5_inp2,F1i2L5_inp3 );

wire F2i2L5_inp1, F2i2L5_inp2, F2i2L5_inp3;
assign F2i2L5_inp1 = sF1i1L5;
assign F2i2L5_inp2 = sF2i1L5;
assign F2i2L5_inp3 = sHi1L5;
wire sF2i2L5, cF2i2L5;
FA F2i2L5( sF2i2L5,cF2i2L5,F2i2L5_inp1,F2i2L5_inp2,F2i2L5_inp3 );

wire F1i2L6_inp1, F1i2L6_inp2, F1i2L6_inp3;
assign F1i2L6_inp1 = cF1i1L5;
assign F1i2L6_inp2 = cF2i1L5;
assign F1i2L6_inp3 = cHi1L5;
wire sF1i2L6, cF1i2L6;
FA F1i2L6( sF1i2L6,cF1i2L6,F1i2L6_inp1,F1i2L6_inp2,F1i2L6_inp3 );

wire F2i2L6_inp1, F2i2L6_inp2, F2i2L6_inp3;
assign F2i2L6_inp1 = sF1i1L6;
assign F2i2L6_inp2 = sF2i1L6;
assign F2i2L6_inp3 = sHi1L6;
wire sF2i2L6, cF2i2L6;
FA F2i2L6( sF2i2L6,cF2i2L6,F2i2L6_inp1,F2i2L6_inp2,F2i2L6_inp3 );

wire F1i2L7_inp1, F1i2L7_inp2, F1i2L7_inp3;
assign F1i2L7_inp1 = cF1i1L6;
assign F1i2L7_inp2 = cF2i1L6;
assign F1i2L7_inp3 = cHi1L6;
wire sF1i2L7, cF1i2L7;
FA F1i2L7( sF1i2L7,cF1i2L7,F1i2L7_inp1,F1i2L7_inp2,F1i2L7_inp3 );

wire F2i2L7_inp1, F2i2L7_inp2, F2i2L7_inp3;
assign F2i2L7_inp1 = sF1i1L7;
assign F2i2L7_inp2 = sF2i1L7;
assign F2i2L7_inp3 = sHi1L7;
wire sF2i2L7, cF2i2L7;
FA F2i2L7( sF2i2L7,cF2i2L7,F2i2L7_inp1,F2i2L7_inp2,F2i2L7_inp3 );

wire F1i2L8_inp1, F1i2L8_inp2, F1i2L8_inp3;
assign F1i2L8_inp1 = cF1i1L7;
assign F1i2L8_inp2 = cF2i1L7;
assign F1i2L8_inp3 = cHi1L7;
wire sF1i2L8, cF1i2L8;
FA F1i2L8( sF1i2L8,cF1i2L8,F1i2L8_inp1,F1i2L8_inp2,F1i2L8_inp3 );

wire F2i2L8_inp1, F2i2L8_inp2, F2i2L8_inp3;
assign F2i2L8_inp1 = sF1i1L8;
assign F2i2L8_inp2 = sF2i1L8;
assign F2i2L8_inp3 = sHi1L8;
wire sF2i2L8, cF2i2L8;
FA F2i2L8( sF2i2L8,cF2i2L8,F2i2L8_inp1,F2i2L8_inp2,F2i2L8_inp3 );

wire F1i2L9_inp1, F1i2L9_inp2, F1i2L9_inp3;
assign F1i2L9_inp1 = cF1i1L8;
assign F1i2L9_inp2 = cF2i1L8;
assign F1i2L9_inp3 = cHi1L8;
wire sF1i2L9, cF1i2L9;
FA F1i2L9( sF1i2L9,cF1i2L9,F1i2L9_inp1,F1i2L9_inp2,F1i2L9_inp3 );

wire F2i2L9_inp1, F2i2L9_inp2, F2i2L9_inp3;
assign F2i2L9_inp1 = sF1i1L9;
assign F2i2L9_inp2 = sF2i1L9;
assign F2i2L9_inp3 = sHi1L9;
wire sF2i2L9, cF2i2L9;
FA F2i2L9( sF2i2L9,cF2i2L9,F2i2L9_inp1,F2i2L9_inp2,F2i2L9_inp3 );

wire F1i2L10_inp1, F1i2L10_inp2, F1i2L10_inp3;
assign F1i2L10_inp1 = cF1i1L9;
assign F1i2L10_inp2 = cF2i1L9;
assign F1i2L10_inp3 = cHi1L9;
wire sF1i2L10, cF1i2L10;
FA F1i2L10( sF1i2L10,cF1i2L10,F1i2L10_inp1,F1i2L10_inp2,F1i2L10_inp3 );

wire F2i2L10_inp1, F2i2L10_inp2, F2i2L10_inp3;
assign F2i2L10_inp1 = sF1i1L10;
assign F2i2L10_inp2 = sF2i1L10;
assign F2i2L10_inp3 = sHi1L10;
wire sF2i2L10, cF2i2L10;
FA F2i2L10( sF2i2L10,cF2i2L10,F2i2L10_inp1,F2i2L10_inp2,F2i2L10_inp3 );

wire F1i2L11_inp1, F1i2L11_inp2, F1i2L11_inp3;
assign F1i2L11_inp1 = cF1i1L10;
assign F1i2L11_inp2 = cF2i1L10;
assign F1i2L11_inp3 = cHi1L10;
wire sF1i2L11, cF1i2L11;
FA F1i2L11( sF1i2L11,cF1i2L11,F1i2L11_inp1,F1i2L11_inp2,F1i2L11_inp3 );

wire F2i2L11_inp1, F2i2L11_inp2, F2i2L11_inp3;
assign F2i2L11_inp1 = sF1i1L11;
assign F2i2L11_inp2 = sF2i1L11;
assign F2i2L11_inp3 = sHi1L11;
wire sF2i2L11, cF2i2L11;
FA F2i2L11( sF2i2L11,cF2i2L11,F2i2L11_inp1,F2i2L11_inp2,F2i2L11_inp3 );

wire Hi2L12_inp1, Hi2L12_inp2;
assign Hi2L12_inp1 = cF1i1L11;
assign Hi2L12_inp2 = cF2i1L11;
wire sHi2L12, cHi2L12;
HA Hi2L12 ( sHi2L12,cHi2L12,Hi2L12_inp1,Hi2L12_inp2 );



///////////// Iteration Number =3///////////////////





wire Hi3L0_inp1, Hi3L0_inp2;
assign Hi3L0_inp1 = G[0];
assign Hi3L0_inp2 = H[0];
wire sHi3L0, cHi3L0;
HA Hi3L0 ( sHi3L0,cHi3L0,Hi3L0_inp1,Hi3L0_inp2 );

wire F1i3L1_inp1, F1i3L1_inp2, F1i3L1_inp3;
assign F1i3L1_inp1 = sHi1L1;
assign F1i3L1_inp2 = cF1i2L0;
assign F1i3L1_inp3 = sF1i2L1;
wire sF1i3L1, cF1i3L1;
FA F1i3L1( sF1i3L1,cF1i3L1,F1i3L1_inp1,F1i3L1_inp2,F1i3L1_inp3 );

wire F1i3L2_inp1, F1i3L2_inp2, F1i3L2_inp3;
assign F1i3L2_inp1 = cF1i2L1;
assign F1i3L2_inp2 = cHi2L1;
assign F1i3L2_inp3 = sF1i2L2;
wire sF1i3L2, cF1i3L2;
FA F1i3L2( sF1i3L2,cF1i3L2,F1i3L2_inp1,F1i3L2_inp2,F1i3L2_inp3 );

wire F1i3L3_inp1, F1i3L3_inp2, F1i3L3_inp3;
assign F1i3L3_inp1 = cF1i2L2;
assign F1i3L3_inp2 = cF2i2L2;
assign F1i3L3_inp3 = sF1i2L3;
wire sF1i3L3, cF1i3L3;
FA F1i3L3( sF1i3L3,cF1i3L3,F1i3L3_inp1,F1i3L3_inp2,F1i3L3_inp3 );

wire F1i3L4_inp1, F1i3L4_inp2, F1i3L4_inp3;
assign F1i3L4_inp1 = cF1i2L3;
assign F1i3L4_inp2 = cF2i2L3;
assign F1i3L4_inp3 = sF1i2L4;
wire sF1i3L4, cF1i3L4;
FA F1i3L4( sF1i3L4,cF1i3L4,F1i3L4_inp1,F1i3L4_inp2,F1i3L4_inp3 );

wire F1i3L5_inp1, F1i3L5_inp2, F1i3L5_inp3;
assign F1i3L5_inp1 = cF1i2L4;
assign F1i3L5_inp2 = cF2i2L4;
assign F1i3L5_inp3 = sF1i2L5;
wire sF1i3L5, cF1i3L5;
FA F1i3L5( sF1i3L5,cF1i3L5,F1i3L5_inp1,F1i3L5_inp2,F1i3L5_inp3 );

wire F1i3L6_inp1, F1i3L6_inp2, F1i3L6_inp3;
assign F1i3L6_inp1 = cF1i2L5;
assign F1i3L6_inp2 = cF2i2L5;
assign F1i3L6_inp3 = sF1i2L6;
wire sF1i3L6, cF1i3L6;
FA F1i3L6( sF1i3L6,cF1i3L6,F1i3L6_inp1,F1i3L6_inp2,F1i3L6_inp3 );

wire F1i3L7_inp1, F1i3L7_inp2, F1i3L7_inp3;
assign F1i3L7_inp1 = cF1i2L6;
assign F1i3L7_inp2 = cF2i2L6;
assign F1i3L7_inp3 = sF1i2L7;
wire sF1i3L7, cF1i3L7;
FA F1i3L7( sF1i3L7,cF1i3L7,F1i3L7_inp1,F1i3L7_inp2,F1i3L7_inp3 );

wire F1i3L8_inp1, F1i3L8_inp2, F1i3L8_inp3;
assign F1i3L8_inp1 = cF1i2L7;
assign F1i3L8_inp2 = cF2i2L7;
assign F1i3L8_inp3 = sF1i2L8;
wire sF1i3L8, cF1i3L8;
FA F1i3L8( sF1i3L8,cF1i3L8,F1i3L8_inp1,F1i3L8_inp2,F1i3L8_inp3 );

wire F1i3L9_inp1, F1i3L9_inp2, F1i3L9_inp3;
assign F1i3L9_inp1 = cF1i2L8;
assign F1i3L9_inp2 = cF2i2L8;
assign F1i3L9_inp3 = sF1i2L9;
wire sF1i3L9, cF1i3L9;
FA F1i3L9( sF1i3L9,cF1i3L9,F1i3L9_inp1,F1i3L9_inp2,F1i3L9_inp3 );

wire F1i3L10_inp1, F1i3L10_inp2, F1i3L10_inp3;
assign F1i3L10_inp1 = cF1i2L9;
assign F1i3L10_inp2 = cF2i2L9;
assign F1i3L10_inp3 = sF1i2L10;
wire sF1i3L10, cF1i3L10;
FA F1i3L10( sF1i3L10,cF1i3L10,F1i3L10_inp1,F1i3L10_inp2,F1i3L10_inp3 );

wire F1i3L11_inp1, F1i3L11_inp2, F1i3L11_inp3;
assign F1i3L11_inp1 = cF1i2L10;
assign F1i3L11_inp2 = cF2i2L10;
assign F1i3L11_inp3 = sF1i2L11;
wire sF1i3L11, cF1i3L11;
FA F1i3L11( sF1i3L11,cF1i3L11,F1i3L11_inp1,F1i3L11_inp2,F1i3L11_inp3 );

wire F1i3L12_inp1, F1i3L12_inp2, F1i3L12_inp3;
assign F1i3L12_inp1 = cHi1L11;
assign F1i3L12_inp2 = cF1i2L11;
assign F1i3L12_inp3 = cF2i2L11;
wire sF1i3L12, cF1i3L12;
FA F1i3L12( sF1i3L12,cF1i3L12,F1i3L12_inp1,F1i3L12_inp2,F1i3L12_inp3 );



///////////// Iteration Number =4///////////////////





wire Hi4L0_inp1, Hi4L0_inp2;
assign Hi4L0_inp1 = sF1i1L0;
assign Hi4L0_inp2 = sF1i2L0;
wire sHi4L0, cHi4L0;
HA Hi4L0 ( sHi4L0,cHi4L0,Hi4L0_inp1,Hi4L0_inp2 );

wire F1i4L1_inp1, F1i4L1_inp2, F1i4L1_inp3;
assign F1i4L1_inp1 = sHi2L1;
assign F1i4L1_inp2 = cHi3L0;
assign F1i4L1_inp3 = sF1i3L1;
wire sF1i4L1, cF1i4L1;
FA F1i4L1( sF1i4L1,cF1i4L1,F1i4L1_inp1,F1i4L1_inp2,F1i4L1_inp3 );

wire F1i4L2_inp1, F1i4L2_inp2, F1i4L2_inp3;
assign F1i4L2_inp1 = sF2i2L2;
assign F1i4L2_inp2 = cF1i3L1;
assign F1i4L2_inp3 = sF1i3L2;
wire sF1i4L2, cF1i4L2;
FA F1i4L2( sF1i4L2,cF1i4L2,F1i4L2_inp1,F1i4L2_inp2,F1i4L2_inp3 );

wire F1i4L3_inp1, F1i4L3_inp2, F1i4L3_inp3;
assign F1i4L3_inp1 = sF2i2L3;
assign F1i4L3_inp2 = cF1i3L2;
assign F1i4L3_inp3 = sF1i3L3;
wire sF1i4L3, cF1i4L3;
FA F1i4L3( sF1i4L3,cF1i4L3,F1i4L3_inp1,F1i4L3_inp2,F1i4L3_inp3 );

wire F1i4L4_inp1, F1i4L4_inp2, F1i4L4_inp3;
assign F1i4L4_inp1 = sF2i2L4;
assign F1i4L4_inp2 = cF1i3L3;
assign F1i4L4_inp3 = sF1i3L4;
wire sF1i4L4, cF1i4L4;
FA F1i4L4( sF1i4L4,cF1i4L4,F1i4L4_inp1,F1i4L4_inp2,F1i4L4_inp3 );

wire F1i4L5_inp1, F1i4L5_inp2, F1i4L5_inp3;
assign F1i4L5_inp1 = sF2i2L5;
assign F1i4L5_inp2 = cF1i3L4;
assign F1i4L5_inp3 = sF1i3L5;
wire sF1i4L5, cF1i4L5;
FA F1i4L5( sF1i4L5,cF1i4L5,F1i4L5_inp1,F1i4L5_inp2,F1i4L5_inp3 );

wire F1i4L6_inp1, F1i4L6_inp2, F1i4L6_inp3;
assign F1i4L6_inp1 = sF2i2L6;
assign F1i4L6_inp2 = cF1i3L5;
assign F1i4L6_inp3 = sF1i3L6;
wire sF1i4L6, cF1i4L6;
FA F1i4L6( sF1i4L6,cF1i4L6,F1i4L6_inp1,F1i4L6_inp2,F1i4L6_inp3 );

wire F1i4L7_inp1, F1i4L7_inp2, F1i4L7_inp3;
assign F1i4L7_inp1 = sF2i2L7;
assign F1i4L7_inp2 = cF1i3L6;
assign F1i4L7_inp3 = sF1i3L7;
wire sF1i4L7, cF1i4L7;
FA F1i4L7( sF1i4L7,cF1i4L7,F1i4L7_inp1,F1i4L7_inp2,F1i4L7_inp3 );

wire F1i4L8_inp1, F1i4L8_inp2, F1i4L8_inp3;
assign F1i4L8_inp1 = sF2i2L8;
assign F1i4L8_inp2 = cF1i3L7;
assign F1i4L8_inp3 = sF1i3L8;
wire sF1i4L8, cF1i4L8;
FA F1i4L8( sF1i4L8,cF1i4L8,F1i4L8_inp1,F1i4L8_inp2,F1i4L8_inp3 );

wire F1i4L9_inp1, F1i4L9_inp2, F1i4L9_inp3;
assign F1i4L9_inp1 = sF2i2L9;
assign F1i4L9_inp2 = cF1i3L8;
assign F1i4L9_inp3 = sF1i3L9;
wire sF1i4L9, cF1i4L9;
FA F1i4L9( sF1i4L9,cF1i4L9,F1i4L9_inp1,F1i4L9_inp2,F1i4L9_inp3 );

wire F1i4L10_inp1, F1i4L10_inp2, F1i4L10_inp3;
assign F1i4L10_inp1 = sF2i2L10;
assign F1i4L10_inp2 = cF1i3L9;
assign F1i4L10_inp3 = sF1i3L10;
wire sF1i4L10, cF1i4L10;
FA F1i4L10( sF1i4L10,cF1i4L10,F1i4L10_inp1,F1i4L10_inp2,F1i4L10_inp3 );

wire F1i4L11_inp1, F1i4L11_inp2, F1i4L11_inp3;
assign F1i4L11_inp1 = sF2i2L11;
assign F1i4L11_inp2 = cF1i3L10;
assign F1i4L11_inp3 = sF1i3L11;
wire sF1i4L11, cF1i4L11;
FA F1i4L11( sF1i4L11,cF1i4L11,F1i4L11_inp1,F1i4L11_inp2,F1i4L11_inp3 );

wire F1i4L12_inp1, F1i4L12_inp2, F1i4L12_inp3;
assign F1i4L12_inp1 = sHi2L12;
assign F1i4L12_inp2 = cF1i3L11;
assign F1i4L12_inp3 = sF1i3L12;
wire sF1i4L12, cF1i4L12;
FA F1i4L12( sF1i4L12,cF1i4L12,F1i4L12_inp1,F1i4L12_inp2,F1i4L12_inp3 );

wire Hi4L13_inp1, Hi4L13_inp2;
assign Hi4L13_inp1 = cHi2L12;
assign Hi4L13_inp2 = cF1i3L12;
wire sHi4L13, cHi4L13;
HA Hi4L13 ( sHi4L13,cHi4L13,Hi4L13_inp1,Hi4L13_inp2 );


assign out1 ={{cHi4L13},{cF1i4L12},{cF1i4L11},{cF1i4L10},{cF1i4L9},{cF1i4L8},{cF1i4L7},{cF1i4L6},{cF1i4L5},{cF1i4L4},{cF1i4L3},{cF1i4L2},{cF1i4L1},{cHi4L0},{sHi3L0}};
assign out2 ={{1'b0},{sHi4L13},{sF1i4L12},{sF1i4L11},{sF1i4L10},{sF1i4L9},{sF1i4L8},{sF1i4L7},{sF1i4L6},{sF1i4L5},{sF1i4L4},{sF1i4L3},{sF1i4L2},{sF1i4L1},{sHi4L0}} ;
endmodule