module adder7x30(
output [32:0] out1,out2,
input [29:0]A,B,C,D,E,F,G );






///////////// Iteration Number =1///////////////////





wire Hi1L0_inp1, Hi1L0_inp2;
assign Hi1L0_inp1 = A[0];
assign Hi1L0_inp2 = B[0];
wire sHi1L0, cHi1L0;
HA Hi1L0 ( sHi1L0,cHi1L0,Hi1L0_inp1,Hi1L0_inp2 );

wire F1i1L1_inp1, F1i1L1_inp2, F1i1L1_inp3;
assign F1i1L1_inp1 = A[1];
assign F1i1L1_inp2 = B[1];
assign F1i1L1_inp3 = C[1];
wire sF1i1L1, cF1i1L1;
FA F1i1L1( sF1i1L1,cF1i1L1,F1i1L1_inp1,F1i1L1_inp2,F1i1L1_inp3 );

wire F1i1L2_inp1, F1i1L2_inp2, F1i1L2_inp3;
assign F1i1L2_inp1 = A[2];
assign F1i1L2_inp2 = B[2];
assign F1i1L2_inp3 = C[2];
wire sF1i1L2, cF1i1L2;
FA F1i1L2( sF1i1L2,cF1i1L2,F1i1L2_inp1,F1i1L2_inp2,F1i1L2_inp3 );

wire F1i1L3_inp1, F1i1L3_inp2, F1i1L3_inp3;
assign F1i1L3_inp1 = A[3];
assign F1i1L3_inp2 = B[3];
assign F1i1L3_inp3 = C[3];
wire sF1i1L3, cF1i1L3;
FA F1i1L3( sF1i1L3,cF1i1L3,F1i1L3_inp1,F1i1L3_inp2,F1i1L3_inp3 );

wire F1i1L4_inp1, F1i1L4_inp2, F1i1L4_inp3;
assign F1i1L4_inp1 = A[4];
assign F1i1L4_inp2 = B[4];
assign F1i1L4_inp3 = C[4];
wire sF1i1L4, cF1i1L4;
FA F1i1L4( sF1i1L4,cF1i1L4,F1i1L4_inp1,F1i1L4_inp2,F1i1L4_inp3 );

wire F1i1L5_inp1, F1i1L5_inp2, F1i1L5_inp3;
assign F1i1L5_inp1 = A[5];
assign F1i1L5_inp2 = B[5];
assign F1i1L5_inp3 = C[5];
wire sF1i1L5, cF1i1L5;
FA F1i1L5( sF1i1L5,cF1i1L5,F1i1L5_inp1,F1i1L5_inp2,F1i1L5_inp3 );

wire F1i1L6_inp1, F1i1L6_inp2, F1i1L6_inp3;
assign F1i1L6_inp1 = A[6];
assign F1i1L6_inp2 = B[6];
assign F1i1L6_inp3 = C[6];
wire sF1i1L6, cF1i1L6;
FA F1i1L6( sF1i1L6,cF1i1L6,F1i1L6_inp1,F1i1L6_inp2,F1i1L6_inp3 );

wire F1i1L7_inp1, F1i1L7_inp2, F1i1L7_inp3;
assign F1i1L7_inp1 = A[7];
assign F1i1L7_inp2 = B[7];
assign F1i1L7_inp3 = C[7];
wire sF1i1L7, cF1i1L7;
FA F1i1L7( sF1i1L7,cF1i1L7,F1i1L7_inp1,F1i1L7_inp2,F1i1L7_inp3 );

wire F1i1L8_inp1, F1i1L8_inp2, F1i1L8_inp3;
assign F1i1L8_inp1 = A[8];
assign F1i1L8_inp2 = B[8];
assign F1i1L8_inp3 = C[8];
wire sF1i1L8, cF1i1L8;
FA F1i1L8( sF1i1L8,cF1i1L8,F1i1L8_inp1,F1i1L8_inp2,F1i1L8_inp3 );

wire F1i1L9_inp1, F1i1L9_inp2, F1i1L9_inp3;
assign F1i1L9_inp1 = A[9];
assign F1i1L9_inp2 = B[9];
assign F1i1L9_inp3 = C[9];
wire sF1i1L9, cF1i1L9;
FA F1i1L9( sF1i1L9,cF1i1L9,F1i1L9_inp1,F1i1L9_inp2,F1i1L9_inp3 );

wire F1i1L10_inp1, F1i1L10_inp2, F1i1L10_inp3;
assign F1i1L10_inp1 = A[10];
assign F1i1L10_inp2 = B[10];
assign F1i1L10_inp3 = C[10];
wire sF1i1L10, cF1i1L10;
FA F1i1L10( sF1i1L10,cF1i1L10,F1i1L10_inp1,F1i1L10_inp2,F1i1L10_inp3 );

wire F1i1L11_inp1, F1i1L11_inp2, F1i1L11_inp3;
assign F1i1L11_inp1 = A[11];
assign F1i1L11_inp2 = B[11];
assign F1i1L11_inp3 = C[11];
wire sF1i1L11, cF1i1L11;
FA F1i1L11( sF1i1L11,cF1i1L11,F1i1L11_inp1,F1i1L11_inp2,F1i1L11_inp3 );

wire F1i1L12_inp1, F1i1L12_inp2, F1i1L12_inp3;
assign F1i1L12_inp1 = A[12];
assign F1i1L12_inp2 = B[12];
assign F1i1L12_inp3 = C[12];
wire sF1i1L12, cF1i1L12;
FA F1i1L12( sF1i1L12,cF1i1L12,F1i1L12_inp1,F1i1L12_inp2,F1i1L12_inp3 );

wire F1i1L13_inp1, F1i1L13_inp2, F1i1L13_inp3;
assign F1i1L13_inp1 = A[13];
assign F1i1L13_inp2 = B[13];
assign F1i1L13_inp3 = C[13];
wire sF1i1L13, cF1i1L13;
FA F1i1L13( sF1i1L13,cF1i1L13,F1i1L13_inp1,F1i1L13_inp2,F1i1L13_inp3 );

wire F1i1L14_inp1, F1i1L14_inp2, F1i1L14_inp3;
assign F1i1L14_inp1 = A[14];
assign F1i1L14_inp2 = B[14];
assign F1i1L14_inp3 = C[14];
wire sF1i1L14, cF1i1L14;
FA F1i1L14( sF1i1L14,cF1i1L14,F1i1L14_inp1,F1i1L14_inp2,F1i1L14_inp3 );

wire F1i1L15_inp1, F1i1L15_inp2, F1i1L15_inp3;
assign F1i1L15_inp1 = A[15];
assign F1i1L15_inp2 = B[15];
assign F1i1L15_inp3 = C[15];
wire sF1i1L15, cF1i1L15;
FA F1i1L15( sF1i1L15,cF1i1L15,F1i1L15_inp1,F1i1L15_inp2,F1i1L15_inp3 );

wire F1i1L16_inp1, F1i1L16_inp2, F1i1L16_inp3;
assign F1i1L16_inp1 = A[16];
assign F1i1L16_inp2 = B[16];
assign F1i1L16_inp3 = C[16];
wire sF1i1L16, cF1i1L16;
FA F1i1L16( sF1i1L16,cF1i1L16,F1i1L16_inp1,F1i1L16_inp2,F1i1L16_inp3 );

wire F1i1L17_inp1, F1i1L17_inp2, F1i1L17_inp3;
assign F1i1L17_inp1 = A[17];
assign F1i1L17_inp2 = B[17];
assign F1i1L17_inp3 = C[17];
wire sF1i1L17, cF1i1L17;
FA F1i1L17( sF1i1L17,cF1i1L17,F1i1L17_inp1,F1i1L17_inp2,F1i1L17_inp3 );

wire F1i1L18_inp1, F1i1L18_inp2, F1i1L18_inp3;
assign F1i1L18_inp1 = A[18];
assign F1i1L18_inp2 = B[18];
assign F1i1L18_inp3 = C[18];
wire sF1i1L18, cF1i1L18;
FA F1i1L18( sF1i1L18,cF1i1L18,F1i1L18_inp1,F1i1L18_inp2,F1i1L18_inp3 );

wire F1i1L19_inp1, F1i1L19_inp2, F1i1L19_inp3;
assign F1i1L19_inp1 = A[19];
assign F1i1L19_inp2 = B[19];
assign F1i1L19_inp3 = C[19];
wire sF1i1L19, cF1i1L19;
FA F1i1L19( sF1i1L19,cF1i1L19,F1i1L19_inp1,F1i1L19_inp2,F1i1L19_inp3 );

wire F1i1L20_inp1, F1i1L20_inp2, F1i1L20_inp3;
assign F1i1L20_inp1 = A[20];
assign F1i1L20_inp2 = B[20];
assign F1i1L20_inp3 = C[20];
wire sF1i1L20, cF1i1L20;
FA F1i1L20( sF1i1L20,cF1i1L20,F1i1L20_inp1,F1i1L20_inp2,F1i1L20_inp3 );

wire F1i1L21_inp1, F1i1L21_inp2, F1i1L21_inp3;
assign F1i1L21_inp1 = A[21];
assign F1i1L21_inp2 = B[21];
assign F1i1L21_inp3 = C[21];
wire sF1i1L21, cF1i1L21;
FA F1i1L21( sF1i1L21,cF1i1L21,F1i1L21_inp1,F1i1L21_inp2,F1i1L21_inp3 );

wire F1i1L22_inp1, F1i1L22_inp2, F1i1L22_inp3;
assign F1i1L22_inp1 = A[22];
assign F1i1L22_inp2 = B[22];
assign F1i1L22_inp3 = C[22];
wire sF1i1L22, cF1i1L22;
FA F1i1L22( sF1i1L22,cF1i1L22,F1i1L22_inp1,F1i1L22_inp2,F1i1L22_inp3 );

wire F1i1L23_inp1, F1i1L23_inp2, F1i1L23_inp3;
assign F1i1L23_inp1 = A[23];
assign F1i1L23_inp2 = B[23];
assign F1i1L23_inp3 = C[23];
wire sF1i1L23, cF1i1L23;
FA F1i1L23( sF1i1L23,cF1i1L23,F1i1L23_inp1,F1i1L23_inp2,F1i1L23_inp3 );

wire F1i1L24_inp1, F1i1L24_inp2, F1i1L24_inp3;
assign F1i1L24_inp1 = A[24];
assign F1i1L24_inp2 = B[24];
assign F1i1L24_inp3 = C[24];
wire sF1i1L24, cF1i1L24;
FA F1i1L24( sF1i1L24,cF1i1L24,F1i1L24_inp1,F1i1L24_inp2,F1i1L24_inp3 );

wire F1i1L25_inp1, F1i1L25_inp2, F1i1L25_inp3;
assign F1i1L25_inp1 = A[25];
assign F1i1L25_inp2 = B[25];
assign F1i1L25_inp3 = C[25];
wire sF1i1L25, cF1i1L25;
FA F1i1L25( sF1i1L25,cF1i1L25,F1i1L25_inp1,F1i1L25_inp2,F1i1L25_inp3 );

wire F1i1L26_inp1, F1i1L26_inp2, F1i1L26_inp3;
assign F1i1L26_inp1 = A[26];
assign F1i1L26_inp2 = B[26];
assign F1i1L26_inp3 = C[26];
wire sF1i1L26, cF1i1L26;
FA F1i1L26( sF1i1L26,cF1i1L26,F1i1L26_inp1,F1i1L26_inp2,F1i1L26_inp3 );

wire F1i1L27_inp1, F1i1L27_inp2, F1i1L27_inp3;
assign F1i1L27_inp1 = A[27];
assign F1i1L27_inp2 = B[27];
assign F1i1L27_inp3 = C[27];
wire sF1i1L27, cF1i1L27;
FA F1i1L27( sF1i1L27,cF1i1L27,F1i1L27_inp1,F1i1L27_inp2,F1i1L27_inp3 );

wire F1i1L28_inp1, F1i1L28_inp2, F1i1L28_inp3;
assign F1i1L28_inp1 = A[28];
assign F1i1L28_inp2 = B[28];
assign F1i1L28_inp3 = C[28];
wire sF1i1L28, cF1i1L28;
FA F1i1L28( sF1i1L28,cF1i1L28,F1i1L28_inp1,F1i1L28_inp2,F1i1L28_inp3 );

wire F1i1L29_inp1, F1i1L29_inp2, F1i1L29_inp3;
assign F1i1L29_inp1 = A[29];
assign F1i1L29_inp2 = B[29];
assign F1i1L29_inp3 = C[29];
wire sF1i1L29, cF1i1L29;
FA F1i1L29( sF1i1L29,cF1i1L29,F1i1L29_inp1,F1i1L29_inp2,F1i1L29_inp3 );



///////////// Iteration Number =2///////////////////





wire F1i2L0_inp1, F1i2L0_inp2, F1i2L0_inp3;
assign F1i2L0_inp1 = C[0];
assign F1i2L0_inp2 = D[0];
assign F1i2L0_inp3 = E[0];
wire sF1i2L0, cF1i2L0;
FA F1i2L0( sF1i2L0,cF1i2L0,F1i2L0_inp1,F1i2L0_inp2,F1i2L0_inp3 );

wire F1i2L1_inp1, F1i2L1_inp2, F1i2L1_inp3;
assign F1i2L1_inp1 = D[1];
assign F1i2L1_inp2 = E[1];
assign F1i2L1_inp3 = F[1];
wire sF1i2L1, cF1i2L1;
FA F1i2L1( sF1i2L1,cF1i2L1,F1i2L1_inp1,F1i2L1_inp2,F1i2L1_inp3 );

wire Hi2L1_inp1, Hi2L1_inp2;
assign Hi2L1_inp1 = G[1];
assign Hi2L1_inp2 = cHi1L0;
wire sHi2L1, cHi2L1;
HA Hi2L1 ( sHi2L1,cHi2L1,Hi2L1_inp1,Hi2L1_inp2 );

wire F1i2L2_inp1, F1i2L2_inp2, F1i2L2_inp3;
assign F1i2L2_inp1 = D[2];
assign F1i2L2_inp2 = E[2];
assign F1i2L2_inp3 = F[2];
wire sF1i2L2, cF1i2L2;
FA F1i2L2( sF1i2L2,cF1i2L2,F1i2L2_inp1,F1i2L2_inp2,F1i2L2_inp3 );

wire F2i2L2_inp1, F2i2L2_inp2, F2i2L2_inp3;
assign F2i2L2_inp1 = G[2];
assign F2i2L2_inp2 = cF1i1L1;
assign F2i2L2_inp3 = sF1i1L2;
wire sF2i2L2, cF2i2L2;
FA F2i2L2( sF2i2L2,cF2i2L2,F2i2L2_inp1,F2i2L2_inp2,F2i2L2_inp3 );

wire F1i2L3_inp1, F1i2L3_inp2, F1i2L3_inp3;
assign F1i2L3_inp1 = D[3];
assign F1i2L3_inp2 = E[3];
assign F1i2L3_inp3 = F[3];
wire sF1i2L3, cF1i2L3;
FA F1i2L3( sF1i2L3,cF1i2L3,F1i2L3_inp1,F1i2L3_inp2,F1i2L3_inp3 );

wire F2i2L3_inp1, F2i2L3_inp2, F2i2L3_inp3;
assign F2i2L3_inp1 = G[3];
assign F2i2L3_inp2 = cF1i1L2;
assign F2i2L3_inp3 = sF1i1L3;
wire sF2i2L3, cF2i2L3;
FA F2i2L3( sF2i2L3,cF2i2L3,F2i2L3_inp1,F2i2L3_inp2,F2i2L3_inp3 );

wire F1i2L4_inp1, F1i2L4_inp2, F1i2L4_inp3;
assign F1i2L4_inp1 = D[4];
assign F1i2L4_inp2 = E[4];
assign F1i2L4_inp3 = F[4];
wire sF1i2L4, cF1i2L4;
FA F1i2L4( sF1i2L4,cF1i2L4,F1i2L4_inp1,F1i2L4_inp2,F1i2L4_inp3 );

wire F2i2L4_inp1, F2i2L4_inp2, F2i2L4_inp3;
assign F2i2L4_inp1 = G[4];
assign F2i2L4_inp2 = cF1i1L3;
assign F2i2L4_inp3 = sF1i1L4;
wire sF2i2L4, cF2i2L4;
FA F2i2L4( sF2i2L4,cF2i2L4,F2i2L4_inp1,F2i2L4_inp2,F2i2L4_inp3 );

wire F1i2L5_inp1, F1i2L5_inp2, F1i2L5_inp3;
assign F1i2L5_inp1 = D[5];
assign F1i2L5_inp2 = E[5];
assign F1i2L5_inp3 = F[5];
wire sF1i2L5, cF1i2L5;
FA F1i2L5( sF1i2L5,cF1i2L5,F1i2L5_inp1,F1i2L5_inp2,F1i2L5_inp3 );

wire F2i2L5_inp1, F2i2L5_inp2, F2i2L5_inp3;
assign F2i2L5_inp1 = G[5];
assign F2i2L5_inp2 = cF1i1L4;
assign F2i2L5_inp3 = sF1i1L5;
wire sF2i2L5, cF2i2L5;
FA F2i2L5( sF2i2L5,cF2i2L5,F2i2L5_inp1,F2i2L5_inp2,F2i2L5_inp3 );

wire F1i2L6_inp1, F1i2L6_inp2, F1i2L6_inp3;
assign F1i2L6_inp1 = D[6];
assign F1i2L6_inp2 = E[6];
assign F1i2L6_inp3 = F[6];
wire sF1i2L6, cF1i2L6;
FA F1i2L6( sF1i2L6,cF1i2L6,F1i2L6_inp1,F1i2L6_inp2,F1i2L6_inp3 );

wire F2i2L6_inp1, F2i2L6_inp2, F2i2L6_inp3;
assign F2i2L6_inp1 = G[6];
assign F2i2L6_inp2 = cF1i1L5;
assign F2i2L6_inp3 = sF1i1L6;
wire sF2i2L6, cF2i2L6;
FA F2i2L6( sF2i2L6,cF2i2L6,F2i2L6_inp1,F2i2L6_inp2,F2i2L6_inp3 );

wire F1i2L7_inp1, F1i2L7_inp2, F1i2L7_inp3;
assign F1i2L7_inp1 = D[7];
assign F1i2L7_inp2 = E[7];
assign F1i2L7_inp3 = F[7];
wire sF1i2L7, cF1i2L7;
FA F1i2L7( sF1i2L7,cF1i2L7,F1i2L7_inp1,F1i2L7_inp2,F1i2L7_inp3 );

wire F2i2L7_inp1, F2i2L7_inp2, F2i2L7_inp3;
assign F2i2L7_inp1 = G[7];
assign F2i2L7_inp2 = cF1i1L6;
assign F2i2L7_inp3 = sF1i1L7;
wire sF2i2L7, cF2i2L7;
FA F2i2L7( sF2i2L7,cF2i2L7,F2i2L7_inp1,F2i2L7_inp2,F2i2L7_inp3 );

wire F1i2L8_inp1, F1i2L8_inp2, F1i2L8_inp3;
assign F1i2L8_inp1 = D[8];
assign F1i2L8_inp2 = E[8];
assign F1i2L8_inp3 = F[8];
wire sF1i2L8, cF1i2L8;
FA F1i2L8( sF1i2L8,cF1i2L8,F1i2L8_inp1,F1i2L8_inp2,F1i2L8_inp3 );

wire F2i2L8_inp1, F2i2L8_inp2, F2i2L8_inp3;
assign F2i2L8_inp1 = G[8];
assign F2i2L8_inp2 = cF1i1L7;
assign F2i2L8_inp3 = sF1i1L8;
wire sF2i2L8, cF2i2L8;
FA F2i2L8( sF2i2L8,cF2i2L8,F2i2L8_inp1,F2i2L8_inp2,F2i2L8_inp3 );

wire F1i2L9_inp1, F1i2L9_inp2, F1i2L9_inp3;
assign F1i2L9_inp1 = D[9];
assign F1i2L9_inp2 = E[9];
assign F1i2L9_inp3 = F[9];
wire sF1i2L9, cF1i2L9;
FA F1i2L9( sF1i2L9,cF1i2L9,F1i2L9_inp1,F1i2L9_inp2,F1i2L9_inp3 );

wire F2i2L9_inp1, F2i2L9_inp2, F2i2L9_inp3;
assign F2i2L9_inp1 = G[9];
assign F2i2L9_inp2 = cF1i1L8;
assign F2i2L9_inp3 = sF1i1L9;
wire sF2i2L9, cF2i2L9;
FA F2i2L9( sF2i2L9,cF2i2L9,F2i2L9_inp1,F2i2L9_inp2,F2i2L9_inp3 );

wire F1i2L10_inp1, F1i2L10_inp2, F1i2L10_inp3;
assign F1i2L10_inp1 = D[10];
assign F1i2L10_inp2 = E[10];
assign F1i2L10_inp3 = F[10];
wire sF1i2L10, cF1i2L10;
FA F1i2L10( sF1i2L10,cF1i2L10,F1i2L10_inp1,F1i2L10_inp2,F1i2L10_inp3 );

wire F2i2L10_inp1, F2i2L10_inp2, F2i2L10_inp3;
assign F2i2L10_inp1 = G[10];
assign F2i2L10_inp2 = cF1i1L9;
assign F2i2L10_inp3 = sF1i1L10;
wire sF2i2L10, cF2i2L10;
FA F2i2L10( sF2i2L10,cF2i2L10,F2i2L10_inp1,F2i2L10_inp2,F2i2L10_inp3 );

wire F1i2L11_inp1, F1i2L11_inp2, F1i2L11_inp3;
assign F1i2L11_inp1 = D[11];
assign F1i2L11_inp2 = E[11];
assign F1i2L11_inp3 = F[11];
wire sF1i2L11, cF1i2L11;
FA F1i2L11( sF1i2L11,cF1i2L11,F1i2L11_inp1,F1i2L11_inp2,F1i2L11_inp3 );

wire F2i2L11_inp1, F2i2L11_inp2, F2i2L11_inp3;
assign F2i2L11_inp1 = G[11];
assign F2i2L11_inp2 = cF1i1L10;
assign F2i2L11_inp3 = sF1i1L11;
wire sF2i2L11, cF2i2L11;
FA F2i2L11( sF2i2L11,cF2i2L11,F2i2L11_inp1,F2i2L11_inp2,F2i2L11_inp3 );

wire F1i2L12_inp1, F1i2L12_inp2, F1i2L12_inp3;
assign F1i2L12_inp1 = D[12];
assign F1i2L12_inp2 = E[12];
assign F1i2L12_inp3 = F[12];
wire sF1i2L12, cF1i2L12;
FA F1i2L12( sF1i2L12,cF1i2L12,F1i2L12_inp1,F1i2L12_inp2,F1i2L12_inp3 );

wire F2i2L12_inp1, F2i2L12_inp2, F2i2L12_inp3;
assign F2i2L12_inp1 = G[12];
assign F2i2L12_inp2 = cF1i1L11;
assign F2i2L12_inp3 = sF1i1L12;
wire sF2i2L12, cF2i2L12;
FA F2i2L12( sF2i2L12,cF2i2L12,F2i2L12_inp1,F2i2L12_inp2,F2i2L12_inp3 );

wire F1i2L13_inp1, F1i2L13_inp2, F1i2L13_inp3;
assign F1i2L13_inp1 = D[13];
assign F1i2L13_inp2 = E[13];
assign F1i2L13_inp3 = F[13];
wire sF1i2L13, cF1i2L13;
FA F1i2L13( sF1i2L13,cF1i2L13,F1i2L13_inp1,F1i2L13_inp2,F1i2L13_inp3 );

wire F2i2L13_inp1, F2i2L13_inp2, F2i2L13_inp3;
assign F2i2L13_inp1 = G[13];
assign F2i2L13_inp2 = cF1i1L12;
assign F2i2L13_inp3 = sF1i1L13;
wire sF2i2L13, cF2i2L13;
FA F2i2L13( sF2i2L13,cF2i2L13,F2i2L13_inp1,F2i2L13_inp2,F2i2L13_inp3 );

wire F1i2L14_inp1, F1i2L14_inp2, F1i2L14_inp3;
assign F1i2L14_inp1 = D[14];
assign F1i2L14_inp2 = E[14];
assign F1i2L14_inp3 = F[14];
wire sF1i2L14, cF1i2L14;
FA F1i2L14( sF1i2L14,cF1i2L14,F1i2L14_inp1,F1i2L14_inp2,F1i2L14_inp3 );

wire F2i2L14_inp1, F2i2L14_inp2, F2i2L14_inp3;
assign F2i2L14_inp1 = G[14];
assign F2i2L14_inp2 = cF1i1L13;
assign F2i2L14_inp3 = sF1i1L14;
wire sF2i2L14, cF2i2L14;
FA F2i2L14( sF2i2L14,cF2i2L14,F2i2L14_inp1,F2i2L14_inp2,F2i2L14_inp3 );

wire F1i2L15_inp1, F1i2L15_inp2, F1i2L15_inp3;
assign F1i2L15_inp1 = D[15];
assign F1i2L15_inp2 = E[15];
assign F1i2L15_inp3 = F[15];
wire sF1i2L15, cF1i2L15;
FA F1i2L15( sF1i2L15,cF1i2L15,F1i2L15_inp1,F1i2L15_inp2,F1i2L15_inp3 );

wire F2i2L15_inp1, F2i2L15_inp2, F2i2L15_inp3;
assign F2i2L15_inp1 = G[15];
assign F2i2L15_inp2 = cF1i1L14;
assign F2i2L15_inp3 = sF1i1L15;
wire sF2i2L15, cF2i2L15;
FA F2i2L15( sF2i2L15,cF2i2L15,F2i2L15_inp1,F2i2L15_inp2,F2i2L15_inp3 );

wire F1i2L16_inp1, F1i2L16_inp2, F1i2L16_inp3;
assign F1i2L16_inp1 = D[16];
assign F1i2L16_inp2 = E[16];
assign F1i2L16_inp3 = F[16];
wire sF1i2L16, cF1i2L16;
FA F1i2L16( sF1i2L16,cF1i2L16,F1i2L16_inp1,F1i2L16_inp2,F1i2L16_inp3 );

wire F2i2L16_inp1, F2i2L16_inp2, F2i2L16_inp3;
assign F2i2L16_inp1 = G[16];
assign F2i2L16_inp2 = cF1i1L15;
assign F2i2L16_inp3 = sF1i1L16;
wire sF2i2L16, cF2i2L16;
FA F2i2L16( sF2i2L16,cF2i2L16,F2i2L16_inp1,F2i2L16_inp2,F2i2L16_inp3 );

wire F1i2L17_inp1, F1i2L17_inp2, F1i2L17_inp3;
assign F1i2L17_inp1 = D[17];
assign F1i2L17_inp2 = E[17];
assign F1i2L17_inp3 = F[17];
wire sF1i2L17, cF1i2L17;
FA F1i2L17( sF1i2L17,cF1i2L17,F1i2L17_inp1,F1i2L17_inp2,F1i2L17_inp3 );

wire F2i2L17_inp1, F2i2L17_inp2, F2i2L17_inp3;
assign F2i2L17_inp1 = G[17];
assign F2i2L17_inp2 = cF1i1L16;
assign F2i2L17_inp3 = sF1i1L17;
wire sF2i2L17, cF2i2L17;
FA F2i2L17( sF2i2L17,cF2i2L17,F2i2L17_inp1,F2i2L17_inp2,F2i2L17_inp3 );

wire F1i2L18_inp1, F1i2L18_inp2, F1i2L18_inp3;
assign F1i2L18_inp1 = D[18];
assign F1i2L18_inp2 = E[18];
assign F1i2L18_inp3 = F[18];
wire sF1i2L18, cF1i2L18;
FA F1i2L18( sF1i2L18,cF1i2L18,F1i2L18_inp1,F1i2L18_inp2,F1i2L18_inp3 );

wire F2i2L18_inp1, F2i2L18_inp2, F2i2L18_inp3;
assign F2i2L18_inp1 = G[18];
assign F2i2L18_inp2 = cF1i1L17;
assign F2i2L18_inp3 = sF1i1L18;
wire sF2i2L18, cF2i2L18;
FA F2i2L18( sF2i2L18,cF2i2L18,F2i2L18_inp1,F2i2L18_inp2,F2i2L18_inp3 );

wire F1i2L19_inp1, F1i2L19_inp2, F1i2L19_inp3;
assign F1i2L19_inp1 = D[19];
assign F1i2L19_inp2 = E[19];
assign F1i2L19_inp3 = F[19];
wire sF1i2L19, cF1i2L19;
FA F1i2L19( sF1i2L19,cF1i2L19,F1i2L19_inp1,F1i2L19_inp2,F1i2L19_inp3 );

wire F2i2L19_inp1, F2i2L19_inp2, F2i2L19_inp3;
assign F2i2L19_inp1 = G[19];
assign F2i2L19_inp2 = cF1i1L18;
assign F2i2L19_inp3 = sF1i1L19;
wire sF2i2L19, cF2i2L19;
FA F2i2L19( sF2i2L19,cF2i2L19,F2i2L19_inp1,F2i2L19_inp2,F2i2L19_inp3 );

wire F1i2L20_inp1, F1i2L20_inp2, F1i2L20_inp3;
assign F1i2L20_inp1 = D[20];
assign F1i2L20_inp2 = E[20];
assign F1i2L20_inp3 = F[20];
wire sF1i2L20, cF1i2L20;
FA F1i2L20( sF1i2L20,cF1i2L20,F1i2L20_inp1,F1i2L20_inp2,F1i2L20_inp3 );

wire F2i2L20_inp1, F2i2L20_inp2, F2i2L20_inp3;
assign F2i2L20_inp1 = G[20];
assign F2i2L20_inp2 = cF1i1L19;
assign F2i2L20_inp3 = sF1i1L20;
wire sF2i2L20, cF2i2L20;
FA F2i2L20( sF2i2L20,cF2i2L20,F2i2L20_inp1,F2i2L20_inp2,F2i2L20_inp3 );

wire F1i2L21_inp1, F1i2L21_inp2, F1i2L21_inp3;
assign F1i2L21_inp1 = D[21];
assign F1i2L21_inp2 = E[21];
assign F1i2L21_inp3 = F[21];
wire sF1i2L21, cF1i2L21;
FA F1i2L21( sF1i2L21,cF1i2L21,F1i2L21_inp1,F1i2L21_inp2,F1i2L21_inp3 );

wire F2i2L21_inp1, F2i2L21_inp2, F2i2L21_inp3;
assign F2i2L21_inp1 = G[21];
assign F2i2L21_inp2 = cF1i1L20;
assign F2i2L21_inp3 = sF1i1L21;
wire sF2i2L21, cF2i2L21;
FA F2i2L21( sF2i2L21,cF2i2L21,F2i2L21_inp1,F2i2L21_inp2,F2i2L21_inp3 );

wire F1i2L22_inp1, F1i2L22_inp2, F1i2L22_inp3;
assign F1i2L22_inp1 = D[22];
assign F1i2L22_inp2 = E[22];
assign F1i2L22_inp3 = F[22];
wire sF1i2L22, cF1i2L22;
FA F1i2L22( sF1i2L22,cF1i2L22,F1i2L22_inp1,F1i2L22_inp2,F1i2L22_inp3 );

wire F2i2L22_inp1, F2i2L22_inp2, F2i2L22_inp3;
assign F2i2L22_inp1 = G[22];
assign F2i2L22_inp2 = cF1i1L21;
assign F2i2L22_inp3 = sF1i1L22;
wire sF2i2L22, cF2i2L22;
FA F2i2L22( sF2i2L22,cF2i2L22,F2i2L22_inp1,F2i2L22_inp2,F2i2L22_inp3 );

wire F1i2L23_inp1, F1i2L23_inp2, F1i2L23_inp3;
assign F1i2L23_inp1 = D[23];
assign F1i2L23_inp2 = E[23];
assign F1i2L23_inp3 = F[23];
wire sF1i2L23, cF1i2L23;
FA F1i2L23( sF1i2L23,cF1i2L23,F1i2L23_inp1,F1i2L23_inp2,F1i2L23_inp3 );

wire F2i2L23_inp1, F2i2L23_inp2, F2i2L23_inp3;
assign F2i2L23_inp1 = G[23];
assign F2i2L23_inp2 = cF1i1L22;
assign F2i2L23_inp3 = sF1i1L23;
wire sF2i2L23, cF2i2L23;
FA F2i2L23( sF2i2L23,cF2i2L23,F2i2L23_inp1,F2i2L23_inp2,F2i2L23_inp3 );

wire F1i2L24_inp1, F1i2L24_inp2, F1i2L24_inp3;
assign F1i2L24_inp1 = D[24];
assign F1i2L24_inp2 = E[24];
assign F1i2L24_inp3 = F[24];
wire sF1i2L24, cF1i2L24;
FA F1i2L24( sF1i2L24,cF1i2L24,F1i2L24_inp1,F1i2L24_inp2,F1i2L24_inp3 );

wire F2i2L24_inp1, F2i2L24_inp2, F2i2L24_inp3;
assign F2i2L24_inp1 = G[24];
assign F2i2L24_inp2 = cF1i1L23;
assign F2i2L24_inp3 = sF1i1L24;
wire sF2i2L24, cF2i2L24;
FA F2i2L24( sF2i2L24,cF2i2L24,F2i2L24_inp1,F2i2L24_inp2,F2i2L24_inp3 );

wire F1i2L25_inp1, F1i2L25_inp2, F1i2L25_inp3;
assign F1i2L25_inp1 = D[25];
assign F1i2L25_inp2 = E[25];
assign F1i2L25_inp3 = F[25];
wire sF1i2L25, cF1i2L25;
FA F1i2L25( sF1i2L25,cF1i2L25,F1i2L25_inp1,F1i2L25_inp2,F1i2L25_inp3 );

wire F2i2L25_inp1, F2i2L25_inp2, F2i2L25_inp3;
assign F2i2L25_inp1 = G[25];
assign F2i2L25_inp2 = cF1i1L24;
assign F2i2L25_inp3 = sF1i1L25;
wire sF2i2L25, cF2i2L25;
FA F2i2L25( sF2i2L25,cF2i2L25,F2i2L25_inp1,F2i2L25_inp2,F2i2L25_inp3 );

wire F1i2L26_inp1, F1i2L26_inp2, F1i2L26_inp3;
assign F1i2L26_inp1 = D[26];
assign F1i2L26_inp2 = E[26];
assign F1i2L26_inp3 = F[26];
wire sF1i2L26, cF1i2L26;
FA F1i2L26( sF1i2L26,cF1i2L26,F1i2L26_inp1,F1i2L26_inp2,F1i2L26_inp3 );

wire F2i2L26_inp1, F2i2L26_inp2, F2i2L26_inp3;
assign F2i2L26_inp1 = G[26];
assign F2i2L26_inp2 = cF1i1L25;
assign F2i2L26_inp3 = sF1i1L26;
wire sF2i2L26, cF2i2L26;
FA F2i2L26( sF2i2L26,cF2i2L26,F2i2L26_inp1,F2i2L26_inp2,F2i2L26_inp3 );

wire F1i2L27_inp1, F1i2L27_inp2, F1i2L27_inp3;
assign F1i2L27_inp1 = D[27];
assign F1i2L27_inp2 = E[27];
assign F1i2L27_inp3 = F[27];
wire sF1i2L27, cF1i2L27;
FA F1i2L27( sF1i2L27,cF1i2L27,F1i2L27_inp1,F1i2L27_inp2,F1i2L27_inp3 );

wire F2i2L27_inp1, F2i2L27_inp2, F2i2L27_inp3;
assign F2i2L27_inp1 = G[27];
assign F2i2L27_inp2 = cF1i1L26;
assign F2i2L27_inp3 = sF1i1L27;
wire sF2i2L27, cF2i2L27;
FA F2i2L27( sF2i2L27,cF2i2L27,F2i2L27_inp1,F2i2L27_inp2,F2i2L27_inp3 );

wire F1i2L28_inp1, F1i2L28_inp2, F1i2L28_inp3;
assign F1i2L28_inp1 = D[28];
assign F1i2L28_inp2 = E[28];
assign F1i2L28_inp3 = F[28];
wire sF1i2L28, cF1i2L28;
FA F1i2L28( sF1i2L28,cF1i2L28,F1i2L28_inp1,F1i2L28_inp2,F1i2L28_inp3 );

wire F2i2L28_inp1, F2i2L28_inp2, F2i2L28_inp3;
assign F2i2L28_inp1 = G[28];
assign F2i2L28_inp2 = cF1i1L27;
assign F2i2L28_inp3 = sF1i1L28;
wire sF2i2L28, cF2i2L28;
FA F2i2L28( sF2i2L28,cF2i2L28,F2i2L28_inp1,F2i2L28_inp2,F2i2L28_inp3 );

wire F1i2L29_inp1, F1i2L29_inp2, F1i2L29_inp3;
assign F1i2L29_inp1 = D[29];
assign F1i2L29_inp2 = E[29];
assign F1i2L29_inp3 = F[29];
wire sF1i2L29, cF1i2L29;
FA F1i2L29( sF1i2L29,cF1i2L29,F1i2L29_inp1,F1i2L29_inp2,F1i2L29_inp3 );

wire F2i2L29_inp1, F2i2L29_inp2, F2i2L29_inp3;
assign F2i2L29_inp1 = G[29];
assign F2i2L29_inp2 = cF1i1L28;
assign F2i2L29_inp3 = sF1i1L29;
wire sF2i2L29, cF2i2L29;
FA F2i2L29( sF2i2L29,cF2i2L29,F2i2L29_inp1,F2i2L29_inp2,F2i2L29_inp3 );



///////////// Iteration Number =3///////////////////





wire Hi3L0_inp1, Hi3L0_inp2;
assign Hi3L0_inp1 = F[0];
assign Hi3L0_inp2 = G[0];
wire sHi3L0, cHi3L0;
HA Hi3L0 ( sHi3L0,cHi3L0,Hi3L0_inp1,Hi3L0_inp2 );

wire F1i3L1_inp1, F1i3L1_inp2, F1i3L1_inp3;
assign F1i3L1_inp1 = sF1i1L1;
assign F1i3L1_inp2 = cF1i2L0;
assign F1i3L1_inp3 = sF1i2L1;
wire sF1i3L1, cF1i3L1;
FA F1i3L1( sF1i3L1,cF1i3L1,F1i3L1_inp1,F1i3L1_inp2,F1i3L1_inp3 );

wire F1i3L2_inp1, F1i3L2_inp2, F1i3L2_inp3;
assign F1i3L2_inp1 = cF1i2L1;
assign F1i3L2_inp2 = cHi2L1;
assign F1i3L2_inp3 = sF1i2L2;
wire sF1i3L2, cF1i3L2;
FA F1i3L2( sF1i3L2,cF1i3L2,F1i3L2_inp1,F1i3L2_inp2,F1i3L2_inp3 );

wire F1i3L3_inp1, F1i3L3_inp2, F1i3L3_inp3;
assign F1i3L3_inp1 = cF1i2L2;
assign F1i3L3_inp2 = cF2i2L2;
assign F1i3L3_inp3 = sF1i2L3;
wire sF1i3L3, cF1i3L3;
FA F1i3L3( sF1i3L3,cF1i3L3,F1i3L3_inp1,F1i3L3_inp2,F1i3L3_inp3 );

wire F1i3L4_inp1, F1i3L4_inp2, F1i3L4_inp3;
assign F1i3L4_inp1 = cF1i2L3;
assign F1i3L4_inp2 = cF2i2L3;
assign F1i3L4_inp3 = sF1i2L4;
wire sF1i3L4, cF1i3L4;
FA F1i3L4( sF1i3L4,cF1i3L4,F1i3L4_inp1,F1i3L4_inp2,F1i3L4_inp3 );

wire F1i3L5_inp1, F1i3L5_inp2, F1i3L5_inp3;
assign F1i3L5_inp1 = cF1i2L4;
assign F1i3L5_inp2 = cF2i2L4;
assign F1i3L5_inp3 = sF1i2L5;
wire sF1i3L5, cF1i3L5;
FA F1i3L5( sF1i3L5,cF1i3L5,F1i3L5_inp1,F1i3L5_inp2,F1i3L5_inp3 );

wire F1i3L6_inp1, F1i3L6_inp2, F1i3L6_inp3;
assign F1i3L6_inp1 = cF1i2L5;
assign F1i3L6_inp2 = cF2i2L5;
assign F1i3L6_inp3 = sF1i2L6;
wire sF1i3L6, cF1i3L6;
FA F1i3L6( sF1i3L6,cF1i3L6,F1i3L6_inp1,F1i3L6_inp2,F1i3L6_inp3 );

wire F1i3L7_inp1, F1i3L7_inp2, F1i3L7_inp3;
assign F1i3L7_inp1 = cF1i2L6;
assign F1i3L7_inp2 = cF2i2L6;
assign F1i3L7_inp3 = sF1i2L7;
wire sF1i3L7, cF1i3L7;
FA F1i3L7( sF1i3L7,cF1i3L7,F1i3L7_inp1,F1i3L7_inp2,F1i3L7_inp3 );

wire F1i3L8_inp1, F1i3L8_inp2, F1i3L8_inp3;
assign F1i3L8_inp1 = cF1i2L7;
assign F1i3L8_inp2 = cF2i2L7;
assign F1i3L8_inp3 = sF1i2L8;
wire sF1i3L8, cF1i3L8;
FA F1i3L8( sF1i3L8,cF1i3L8,F1i3L8_inp1,F1i3L8_inp2,F1i3L8_inp3 );

wire F1i3L9_inp1, F1i3L9_inp2, F1i3L9_inp3;
assign F1i3L9_inp1 = cF1i2L8;
assign F1i3L9_inp2 = cF2i2L8;
assign F1i3L9_inp3 = sF1i2L9;
wire sF1i3L9, cF1i3L9;
FA F1i3L9( sF1i3L9,cF1i3L9,F1i3L9_inp1,F1i3L9_inp2,F1i3L9_inp3 );

wire F1i3L10_inp1, F1i3L10_inp2, F1i3L10_inp3;
assign F1i3L10_inp1 = cF1i2L9;
assign F1i3L10_inp2 = cF2i2L9;
assign F1i3L10_inp3 = sF1i2L10;
wire sF1i3L10, cF1i3L10;
FA F1i3L10( sF1i3L10,cF1i3L10,F1i3L10_inp1,F1i3L10_inp2,F1i3L10_inp3 );

wire F1i3L11_inp1, F1i3L11_inp2, F1i3L11_inp3;
assign F1i3L11_inp1 = cF1i2L10;
assign F1i3L11_inp2 = cF2i2L10;
assign F1i3L11_inp3 = sF1i2L11;
wire sF1i3L11, cF1i3L11;
FA F1i3L11( sF1i3L11,cF1i3L11,F1i3L11_inp1,F1i3L11_inp2,F1i3L11_inp3 );

wire F1i3L12_inp1, F1i3L12_inp2, F1i3L12_inp3;
assign F1i3L12_inp1 = cF1i2L11;
assign F1i3L12_inp2 = cF2i2L11;
assign F1i3L12_inp3 = sF1i2L12;
wire sF1i3L12, cF1i3L12;
FA F1i3L12( sF1i3L12,cF1i3L12,F1i3L12_inp1,F1i3L12_inp2,F1i3L12_inp3 );

wire F1i3L13_inp1, F1i3L13_inp2, F1i3L13_inp3;
assign F1i3L13_inp1 = cF1i2L12;
assign F1i3L13_inp2 = cF2i2L12;
assign F1i3L13_inp3 = sF1i2L13;
wire sF1i3L13, cF1i3L13;
FA F1i3L13( sF1i3L13,cF1i3L13,F1i3L13_inp1,F1i3L13_inp2,F1i3L13_inp3 );

wire F1i3L14_inp1, F1i3L14_inp2, F1i3L14_inp3;
assign F1i3L14_inp1 = cF1i2L13;
assign F1i3L14_inp2 = cF2i2L13;
assign F1i3L14_inp3 = sF1i2L14;
wire sF1i3L14, cF1i3L14;
FA F1i3L14( sF1i3L14,cF1i3L14,F1i3L14_inp1,F1i3L14_inp2,F1i3L14_inp3 );

wire F1i3L15_inp1, F1i3L15_inp2, F1i3L15_inp3;
assign F1i3L15_inp1 = cF1i2L14;
assign F1i3L15_inp2 = cF2i2L14;
assign F1i3L15_inp3 = sF1i2L15;
wire sF1i3L15, cF1i3L15;
FA F1i3L15( sF1i3L15,cF1i3L15,F1i3L15_inp1,F1i3L15_inp2,F1i3L15_inp3 );

wire F1i3L16_inp1, F1i3L16_inp2, F1i3L16_inp3;
assign F1i3L16_inp1 = cF1i2L15;
assign F1i3L16_inp2 = cF2i2L15;
assign F1i3L16_inp3 = sF1i2L16;
wire sF1i3L16, cF1i3L16;
FA F1i3L16( sF1i3L16,cF1i3L16,F1i3L16_inp1,F1i3L16_inp2,F1i3L16_inp3 );

wire F1i3L17_inp1, F1i3L17_inp2, F1i3L17_inp3;
assign F1i3L17_inp1 = cF1i2L16;
assign F1i3L17_inp2 = cF2i2L16;
assign F1i3L17_inp3 = sF1i2L17;
wire sF1i3L17, cF1i3L17;
FA F1i3L17( sF1i3L17,cF1i3L17,F1i3L17_inp1,F1i3L17_inp2,F1i3L17_inp3 );

wire F1i3L18_inp1, F1i3L18_inp2, F1i3L18_inp3;
assign F1i3L18_inp1 = cF1i2L17;
assign F1i3L18_inp2 = cF2i2L17;
assign F1i3L18_inp3 = sF1i2L18;
wire sF1i3L18, cF1i3L18;
FA F1i3L18( sF1i3L18,cF1i3L18,F1i3L18_inp1,F1i3L18_inp2,F1i3L18_inp3 );

wire F1i3L19_inp1, F1i3L19_inp2, F1i3L19_inp3;
assign F1i3L19_inp1 = cF1i2L18;
assign F1i3L19_inp2 = cF2i2L18;
assign F1i3L19_inp3 = sF1i2L19;
wire sF1i3L19, cF1i3L19;
FA F1i3L19( sF1i3L19,cF1i3L19,F1i3L19_inp1,F1i3L19_inp2,F1i3L19_inp3 );

wire F1i3L20_inp1, F1i3L20_inp2, F1i3L20_inp3;
assign F1i3L20_inp1 = cF1i2L19;
assign F1i3L20_inp2 = cF2i2L19;
assign F1i3L20_inp3 = sF1i2L20;
wire sF1i3L20, cF1i3L20;
FA F1i3L20( sF1i3L20,cF1i3L20,F1i3L20_inp1,F1i3L20_inp2,F1i3L20_inp3 );

wire F1i3L21_inp1, F1i3L21_inp2, F1i3L21_inp3;
assign F1i3L21_inp1 = cF1i2L20;
assign F1i3L21_inp2 = cF2i2L20;
assign F1i3L21_inp3 = sF1i2L21;
wire sF1i3L21, cF1i3L21;
FA F1i3L21( sF1i3L21,cF1i3L21,F1i3L21_inp1,F1i3L21_inp2,F1i3L21_inp3 );

wire F1i3L22_inp1, F1i3L22_inp2, F1i3L22_inp3;
assign F1i3L22_inp1 = cF1i2L21;
assign F1i3L22_inp2 = cF2i2L21;
assign F1i3L22_inp3 = sF1i2L22;
wire sF1i3L22, cF1i3L22;
FA F1i3L22( sF1i3L22,cF1i3L22,F1i3L22_inp1,F1i3L22_inp2,F1i3L22_inp3 );

wire F1i3L23_inp1, F1i3L23_inp2, F1i3L23_inp3;
assign F1i3L23_inp1 = cF1i2L22;
assign F1i3L23_inp2 = cF2i2L22;
assign F1i3L23_inp3 = sF1i2L23;
wire sF1i3L23, cF1i3L23;
FA F1i3L23( sF1i3L23,cF1i3L23,F1i3L23_inp1,F1i3L23_inp2,F1i3L23_inp3 );

wire F1i3L24_inp1, F1i3L24_inp2, F1i3L24_inp3;
assign F1i3L24_inp1 = cF1i2L23;
assign F1i3L24_inp2 = cF2i2L23;
assign F1i3L24_inp3 = sF1i2L24;
wire sF1i3L24, cF1i3L24;
FA F1i3L24( sF1i3L24,cF1i3L24,F1i3L24_inp1,F1i3L24_inp2,F1i3L24_inp3 );

wire F1i3L25_inp1, F1i3L25_inp2, F1i3L25_inp3;
assign F1i3L25_inp1 = cF1i2L24;
assign F1i3L25_inp2 = cF2i2L24;
assign F1i3L25_inp3 = sF1i2L25;
wire sF1i3L25, cF1i3L25;
FA F1i3L25( sF1i3L25,cF1i3L25,F1i3L25_inp1,F1i3L25_inp2,F1i3L25_inp3 );

wire F1i3L26_inp1, F1i3L26_inp2, F1i3L26_inp3;
assign F1i3L26_inp1 = cF1i2L25;
assign F1i3L26_inp2 = cF2i2L25;
assign F1i3L26_inp3 = sF1i2L26;
wire sF1i3L26, cF1i3L26;
FA F1i3L26( sF1i3L26,cF1i3L26,F1i3L26_inp1,F1i3L26_inp2,F1i3L26_inp3 );

wire F1i3L27_inp1, F1i3L27_inp2, F1i3L27_inp3;
assign F1i3L27_inp1 = cF1i2L26;
assign F1i3L27_inp2 = cF2i2L26;
assign F1i3L27_inp3 = sF1i2L27;
wire sF1i3L27, cF1i3L27;
FA F1i3L27( sF1i3L27,cF1i3L27,F1i3L27_inp1,F1i3L27_inp2,F1i3L27_inp3 );

wire F1i3L28_inp1, F1i3L28_inp2, F1i3L28_inp3;
assign F1i3L28_inp1 = cF1i2L27;
assign F1i3L28_inp2 = cF2i2L27;
assign F1i3L28_inp3 = sF1i2L28;
wire sF1i3L28, cF1i3L28;
FA F1i3L28( sF1i3L28,cF1i3L28,F1i3L28_inp1,F1i3L28_inp2,F1i3L28_inp3 );

wire F1i3L29_inp1, F1i3L29_inp2, F1i3L29_inp3;
assign F1i3L29_inp1 = cF1i2L28;
assign F1i3L29_inp2 = cF2i2L28;
assign F1i3L29_inp3 = sF1i2L29;
wire sF1i3L29, cF1i3L29;
FA F1i3L29( sF1i3L29,cF1i3L29,F1i3L29_inp1,F1i3L29_inp2,F1i3L29_inp3 );

wire Hi3L30_inp1, Hi3L30_inp2;
assign Hi3L30_inp1 = cF1i1L29;
assign Hi3L30_inp2 = cF1i2L29;
wire sHi3L30, cHi3L30;
HA Hi3L30 ( sHi3L30,cHi3L30,Hi3L30_inp1,Hi3L30_inp2 );



///////////// Iteration Number =4///////////////////





wire Hi4L0_inp1, Hi4L0_inp2;
assign Hi4L0_inp1 = sHi1L0;
assign Hi4L0_inp2 = sF1i2L0;
wire sHi4L0, cHi4L0;
HA Hi4L0 ( sHi4L0,cHi4L0,Hi4L0_inp1,Hi4L0_inp2 );

wire F1i4L1_inp1, F1i4L1_inp2, F1i4L1_inp3;
assign F1i4L1_inp1 = sHi2L1;
assign F1i4L1_inp2 = cHi3L0;
assign F1i4L1_inp3 = sF1i3L1;
wire sF1i4L1, cF1i4L1;
FA F1i4L1( sF1i4L1,cF1i4L1,F1i4L1_inp1,F1i4L1_inp2,F1i4L1_inp3 );

wire F1i4L2_inp1, F1i4L2_inp2, F1i4L2_inp3;
assign F1i4L2_inp1 = sF2i2L2;
assign F1i4L2_inp2 = cF1i3L1;
assign F1i4L2_inp3 = sF1i3L2;
wire sF1i4L2, cF1i4L2;
FA F1i4L2( sF1i4L2,cF1i4L2,F1i4L2_inp1,F1i4L2_inp2,F1i4L2_inp3 );

wire F1i4L3_inp1, F1i4L3_inp2, F1i4L3_inp3;
assign F1i4L3_inp1 = sF2i2L3;
assign F1i4L3_inp2 = cF1i3L2;
assign F1i4L3_inp3 = sF1i3L3;
wire sF1i4L3, cF1i4L3;
FA F1i4L3( sF1i4L3,cF1i4L3,F1i4L3_inp1,F1i4L3_inp2,F1i4L3_inp3 );

wire F1i4L4_inp1, F1i4L4_inp2, F1i4L4_inp3;
assign F1i4L4_inp1 = sF2i2L4;
assign F1i4L4_inp2 = cF1i3L3;
assign F1i4L4_inp3 = sF1i3L4;
wire sF1i4L4, cF1i4L4;
FA F1i4L4( sF1i4L4,cF1i4L4,F1i4L4_inp1,F1i4L4_inp2,F1i4L4_inp3 );

wire F1i4L5_inp1, F1i4L5_inp2, F1i4L5_inp3;
assign F1i4L5_inp1 = sF2i2L5;
assign F1i4L5_inp2 = cF1i3L4;
assign F1i4L5_inp3 = sF1i3L5;
wire sF1i4L5, cF1i4L5;
FA F1i4L5( sF1i4L5,cF1i4L5,F1i4L5_inp1,F1i4L5_inp2,F1i4L5_inp3 );

wire F1i4L6_inp1, F1i4L6_inp2, F1i4L6_inp3;
assign F1i4L6_inp1 = sF2i2L6;
assign F1i4L6_inp2 = cF1i3L5;
assign F1i4L6_inp3 = sF1i3L6;
wire sF1i4L6, cF1i4L6;
FA F1i4L6( sF1i4L6,cF1i4L6,F1i4L6_inp1,F1i4L6_inp2,F1i4L6_inp3 );

wire F1i4L7_inp1, F1i4L7_inp2, F1i4L7_inp3;
assign F1i4L7_inp1 = sF2i2L7;
assign F1i4L7_inp2 = cF1i3L6;
assign F1i4L7_inp3 = sF1i3L7;
wire sF1i4L7, cF1i4L7;
FA F1i4L7( sF1i4L7,cF1i4L7,F1i4L7_inp1,F1i4L7_inp2,F1i4L7_inp3 );

wire F1i4L8_inp1, F1i4L8_inp2, F1i4L8_inp3;
assign F1i4L8_inp1 = sF2i2L8;
assign F1i4L8_inp2 = cF1i3L7;
assign F1i4L8_inp3 = sF1i3L8;
wire sF1i4L8, cF1i4L8;
FA F1i4L8( sF1i4L8,cF1i4L8,F1i4L8_inp1,F1i4L8_inp2,F1i4L8_inp3 );

wire F1i4L9_inp1, F1i4L9_inp2, F1i4L9_inp3;
assign F1i4L9_inp1 = sF2i2L9;
assign F1i4L9_inp2 = cF1i3L8;
assign F1i4L9_inp3 = sF1i3L9;
wire sF1i4L9, cF1i4L9;
FA F1i4L9( sF1i4L9,cF1i4L9,F1i4L9_inp1,F1i4L9_inp2,F1i4L9_inp3 );

wire F1i4L10_inp1, F1i4L10_inp2, F1i4L10_inp3;
assign F1i4L10_inp1 = sF2i2L10;
assign F1i4L10_inp2 = cF1i3L9;
assign F1i4L10_inp3 = sF1i3L10;
wire sF1i4L10, cF1i4L10;
FA F1i4L10( sF1i4L10,cF1i4L10,F1i4L10_inp1,F1i4L10_inp2,F1i4L10_inp3 );

wire F1i4L11_inp1, F1i4L11_inp2, F1i4L11_inp3;
assign F1i4L11_inp1 = sF2i2L11;
assign F1i4L11_inp2 = cF1i3L10;
assign F1i4L11_inp3 = sF1i3L11;
wire sF1i4L11, cF1i4L11;
FA F1i4L11( sF1i4L11,cF1i4L11,F1i4L11_inp1,F1i4L11_inp2,F1i4L11_inp3 );

wire F1i4L12_inp1, F1i4L12_inp2, F1i4L12_inp3;
assign F1i4L12_inp1 = sF2i2L12;
assign F1i4L12_inp2 = cF1i3L11;
assign F1i4L12_inp3 = sF1i3L12;
wire sF1i4L12, cF1i4L12;
FA F1i4L12( sF1i4L12,cF1i4L12,F1i4L12_inp1,F1i4L12_inp2,F1i4L12_inp3 );

wire F1i4L13_inp1, F1i4L13_inp2, F1i4L13_inp3;
assign F1i4L13_inp1 = sF2i2L13;
assign F1i4L13_inp2 = cF1i3L12;
assign F1i4L13_inp3 = sF1i3L13;
wire sF1i4L13, cF1i4L13;
FA F1i4L13( sF1i4L13,cF1i4L13,F1i4L13_inp1,F1i4L13_inp2,F1i4L13_inp3 );

wire F1i4L14_inp1, F1i4L14_inp2, F1i4L14_inp3;
assign F1i4L14_inp1 = sF2i2L14;
assign F1i4L14_inp2 = cF1i3L13;
assign F1i4L14_inp3 = sF1i3L14;
wire sF1i4L14, cF1i4L14;
FA F1i4L14( sF1i4L14,cF1i4L14,F1i4L14_inp1,F1i4L14_inp2,F1i4L14_inp3 );

wire F1i4L15_inp1, F1i4L15_inp2, F1i4L15_inp3;
assign F1i4L15_inp1 = sF2i2L15;
assign F1i4L15_inp2 = cF1i3L14;
assign F1i4L15_inp3 = sF1i3L15;
wire sF1i4L15, cF1i4L15;
FA F1i4L15( sF1i4L15,cF1i4L15,F1i4L15_inp1,F1i4L15_inp2,F1i4L15_inp3 );

wire F1i4L16_inp1, F1i4L16_inp2, F1i4L16_inp3;
assign F1i4L16_inp1 = sF2i2L16;
assign F1i4L16_inp2 = cF1i3L15;
assign F1i4L16_inp3 = sF1i3L16;
wire sF1i4L16, cF1i4L16;
FA F1i4L16( sF1i4L16,cF1i4L16,F1i4L16_inp1,F1i4L16_inp2,F1i4L16_inp3 );

wire F1i4L17_inp1, F1i4L17_inp2, F1i4L17_inp3;
assign F1i4L17_inp1 = sF2i2L17;
assign F1i4L17_inp2 = cF1i3L16;
assign F1i4L17_inp3 = sF1i3L17;
wire sF1i4L17, cF1i4L17;
FA F1i4L17( sF1i4L17,cF1i4L17,F1i4L17_inp1,F1i4L17_inp2,F1i4L17_inp3 );

wire F1i4L18_inp1, F1i4L18_inp2, F1i4L18_inp3;
assign F1i4L18_inp1 = sF2i2L18;
assign F1i4L18_inp2 = cF1i3L17;
assign F1i4L18_inp3 = sF1i3L18;
wire sF1i4L18, cF1i4L18;
FA F1i4L18( sF1i4L18,cF1i4L18,F1i4L18_inp1,F1i4L18_inp2,F1i4L18_inp3 );

wire F1i4L19_inp1, F1i4L19_inp2, F1i4L19_inp3;
assign F1i4L19_inp1 = sF2i2L19;
assign F1i4L19_inp2 = cF1i3L18;
assign F1i4L19_inp3 = sF1i3L19;
wire sF1i4L19, cF1i4L19;
FA F1i4L19( sF1i4L19,cF1i4L19,F1i4L19_inp1,F1i4L19_inp2,F1i4L19_inp3 );

wire F1i4L20_inp1, F1i4L20_inp2, F1i4L20_inp3;
assign F1i4L20_inp1 = sF2i2L20;
assign F1i4L20_inp2 = cF1i3L19;
assign F1i4L20_inp3 = sF1i3L20;
wire sF1i4L20, cF1i4L20;
FA F1i4L20( sF1i4L20,cF1i4L20,F1i4L20_inp1,F1i4L20_inp2,F1i4L20_inp3 );

wire F1i4L21_inp1, F1i4L21_inp2, F1i4L21_inp3;
assign F1i4L21_inp1 = sF2i2L21;
assign F1i4L21_inp2 = cF1i3L20;
assign F1i4L21_inp3 = sF1i3L21;
wire sF1i4L21, cF1i4L21;
FA F1i4L21( sF1i4L21,cF1i4L21,F1i4L21_inp1,F1i4L21_inp2,F1i4L21_inp3 );

wire F1i4L22_inp1, F1i4L22_inp2, F1i4L22_inp3;
assign F1i4L22_inp1 = sF2i2L22;
assign F1i4L22_inp2 = cF1i3L21;
assign F1i4L22_inp3 = sF1i3L22;
wire sF1i4L22, cF1i4L22;
FA F1i4L22( sF1i4L22,cF1i4L22,F1i4L22_inp1,F1i4L22_inp2,F1i4L22_inp3 );

wire F1i4L23_inp1, F1i4L23_inp2, F1i4L23_inp3;
assign F1i4L23_inp1 = sF2i2L23;
assign F1i4L23_inp2 = cF1i3L22;
assign F1i4L23_inp3 = sF1i3L23;
wire sF1i4L23, cF1i4L23;
FA F1i4L23( sF1i4L23,cF1i4L23,F1i4L23_inp1,F1i4L23_inp2,F1i4L23_inp3 );

wire F1i4L24_inp1, F1i4L24_inp2, F1i4L24_inp3;
assign F1i4L24_inp1 = sF2i2L24;
assign F1i4L24_inp2 = cF1i3L23;
assign F1i4L24_inp3 = sF1i3L24;
wire sF1i4L24, cF1i4L24;
FA F1i4L24( sF1i4L24,cF1i4L24,F1i4L24_inp1,F1i4L24_inp2,F1i4L24_inp3 );

wire F1i4L25_inp1, F1i4L25_inp2, F1i4L25_inp3;
assign F1i4L25_inp1 = sF2i2L25;
assign F1i4L25_inp2 = cF1i3L24;
assign F1i4L25_inp3 = sF1i3L25;
wire sF1i4L25, cF1i4L25;
FA F1i4L25( sF1i4L25,cF1i4L25,F1i4L25_inp1,F1i4L25_inp2,F1i4L25_inp3 );

wire F1i4L26_inp1, F1i4L26_inp2, F1i4L26_inp3;
assign F1i4L26_inp1 = sF2i2L26;
assign F1i4L26_inp2 = cF1i3L25;
assign F1i4L26_inp3 = sF1i3L26;
wire sF1i4L26, cF1i4L26;
FA F1i4L26( sF1i4L26,cF1i4L26,F1i4L26_inp1,F1i4L26_inp2,F1i4L26_inp3 );

wire F1i4L27_inp1, F1i4L27_inp2, F1i4L27_inp3;
assign F1i4L27_inp1 = sF2i2L27;
assign F1i4L27_inp2 = cF1i3L26;
assign F1i4L27_inp3 = sF1i3L27;
wire sF1i4L27, cF1i4L27;
FA F1i4L27( sF1i4L27,cF1i4L27,F1i4L27_inp1,F1i4L27_inp2,F1i4L27_inp3 );

wire F1i4L28_inp1, F1i4L28_inp2, F1i4L28_inp3;
assign F1i4L28_inp1 = sF2i2L28;
assign F1i4L28_inp2 = cF1i3L27;
assign F1i4L28_inp3 = sF1i3L28;
wire sF1i4L28, cF1i4L28;
FA F1i4L28( sF1i4L28,cF1i4L28,F1i4L28_inp1,F1i4L28_inp2,F1i4L28_inp3 );

wire F1i4L29_inp1, F1i4L29_inp2, F1i4L29_inp3;
assign F1i4L29_inp1 = sF2i2L29;
assign F1i4L29_inp2 = cF1i3L28;
assign F1i4L29_inp3 = sF1i3L29;
wire sF1i4L29, cF1i4L29;
FA F1i4L29( sF1i4L29,cF1i4L29,F1i4L29_inp1,F1i4L29_inp2,F1i4L29_inp3 );

wire F1i4L30_inp1, F1i4L30_inp2, F1i4L30_inp3;
assign F1i4L30_inp1 = cF2i2L29;
assign F1i4L30_inp2 = cF1i3L29;
assign F1i4L30_inp3 = sHi3L30;
wire sF1i4L30, cF1i4L30;
FA F1i4L30( sF1i4L30,cF1i4L30,F1i4L30_inp1,F1i4L30_inp2,F1i4L30_inp3 );


assign out1 ={{1'b0},{cHi3L30},{cF1i4L29},{cF1i4L28},{cF1i4L27},{cF1i4L26},{cF1i4L25},{cF1i4L24},{cF1i4L23},{cF1i4L22},{cF1i4L21},{cF1i4L20},{cF1i4L19},{cF1i4L18},{cF1i4L17},{cF1i4L16},{cF1i4L15},{cF1i4L14},{cF1i4L13},{cF1i4L12},{cF1i4L11},{cF1i4L10},{cF1i4L9},{cF1i4L8},{cF1i4L7},{cF1i4L6},{cF1i4L5},{cF1i4L4},{cF1i4L3},{cF1i4L2},{cF1i4L1},{cHi4L0},{sHi3L0}};
assign out2 ={{1'b0},{cF1i4L30},{sF1i4L30},{sF1i4L29},{sF1i4L28},{sF1i4L27},{sF1i4L26},{sF1i4L25},{sF1i4L24},{sF1i4L23},{sF1i4L22},{sF1i4L21},{sF1i4L20},{sF1i4L19},{sF1i4L18},{sF1i4L17},{sF1i4L16},{sF1i4L15},{sF1i4L14},{sF1i4L13},{sF1i4L12},{sF1i4L11},{sF1i4L10},{sF1i4L9},{sF1i4L8},{sF1i4L7},{sF1i4L6},{sF1i4L5},{sF1i4L4},{sF1i4L3},{sF1i4L2},{sF1i4L1},{sHi4L0}} ;
endmodule