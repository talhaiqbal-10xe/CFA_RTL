module mult14x16(
output [29:0] out1,out2,
input [13:0] A,
input [15:0] B );


wire [29:0] CV;
 assign CV=30'b100000000000000010000000000000;
integer i;
 reg[13:0] PP[ 0:15];
always@*
begin
   for ( i=0 ; i<16; i = i+1 )
   begin
      PP[i]= A & {14{B[i]}};
   end
end



///////////// Iteration Number =1///////////////////





wire F1i1L13_inp1, F1i1L13_inp2, F1i1L13_inp3;
assign F1i1L13_inp1 = ~PP[0][13];
assign F1i1L13_inp2 = PP[1][12];
assign F1i1L13_inp3 = PP[2][11];
wire sF1i1L13, cF1i1L13;
FA F1i1L13( sF1i1L13,cF1i1L13,F1i1L13_inp1,F1i1L13_inp2,F1i1L13_inp3 );

wire F1i1L14_inp1, F1i1L14_inp2, F1i1L14_inp3;
assign F1i1L14_inp1 = ~PP[1][13];
assign F1i1L14_inp2 = PP[2][12];
assign F1i1L14_inp3 = PP[3][11];
wire sF1i1L14, cF1i1L14;
FA F1i1L14( sF1i1L14,cF1i1L14,F1i1L14_inp1,F1i1L14_inp2,F1i1L14_inp3 );

wire F1i1L15_inp1, F1i1L15_inp2, F1i1L15_inp3;
assign F1i1L15_inp1 = ~PP[2][13];
assign F1i1L15_inp2 = PP[3][12];
assign F1i1L15_inp3 = PP[4][11];
wire sF1i1L15, cF1i1L15;
FA F1i1L15( sF1i1L15,cF1i1L15,F1i1L15_inp1,F1i1L15_inp2,F1i1L15_inp3 );

wire Hi1L16_inp1, Hi1L16_inp2;
assign Hi1L16_inp1 = ~PP[3][13];
assign Hi1L16_inp2 = PP[4][12];
wire sHi1L16, cHi1L16;
HA Hi1L16 ( sHi1L16,cHi1L16,Hi1L16_inp1,Hi1L16_inp2 );



///////////// Iteration Number =2///////////////////





wire Hi2L9_inp1, Hi2L9_inp2;
assign Hi2L9_inp1 = PP[0][9];
assign Hi2L9_inp2 = PP[1][8];
wire sHi2L9, cHi2L9;
HA Hi2L9 ( sHi2L9,cHi2L9,Hi2L9_inp1,Hi2L9_inp2 );

wire F1i2L10_inp1, F1i2L10_inp2, F1i2L10_inp3;
assign F1i2L10_inp1 = PP[0][10];
assign F1i2L10_inp2 = PP[1][9];
assign F1i2L10_inp3 = PP[2][8];
wire sF1i2L10, cF1i2L10;
FA F1i2L10( sF1i2L10,cF1i2L10,F1i2L10_inp1,F1i2L10_inp2,F1i2L10_inp3 );

wire Hi2L10_inp1, Hi2L10_inp2;
assign Hi2L10_inp1 = PP[3][7];
assign Hi2L10_inp2 = PP[4][6];
wire sHi2L10, cHi2L10;
HA Hi2L10 ( sHi2L10,cHi2L10,Hi2L10_inp1,Hi2L10_inp2 );

wire F1i2L11_inp1, F1i2L11_inp2, F1i2L11_inp3;
assign F1i2L11_inp1 = PP[0][11];
assign F1i2L11_inp2 = PP[1][10];
assign F1i2L11_inp3 = PP[2][9];
wire sF1i2L11, cF1i2L11;
FA F1i2L11( sF1i2L11,cF1i2L11,F1i2L11_inp1,F1i2L11_inp2,F1i2L11_inp3 );

wire F2i2L11_inp1, F2i2L11_inp2, F2i2L11_inp3;
assign F2i2L11_inp1 = PP[3][8];
assign F2i2L11_inp2 = PP[4][7];
assign F2i2L11_inp3 = PP[5][6];
wire sF2i2L11, cF2i2L11;
FA F2i2L11( sF2i2L11,cF2i2L11,F2i2L11_inp1,F2i2L11_inp2,F2i2L11_inp3 );

wire Hi2L11_inp1, Hi2L11_inp2;
assign Hi2L11_inp1 = PP[6][5];
assign Hi2L11_inp2 = PP[7][4];
wire sHi2L11, cHi2L11;
HA Hi2L11 ( sHi2L11,cHi2L11,Hi2L11_inp1,Hi2L11_inp2 );

wire F1i2L12_inp1, F1i2L12_inp2, F1i2L12_inp3;
assign F1i2L12_inp1 = PP[0][12];
assign F1i2L12_inp2 = PP[1][11];
assign F1i2L12_inp3 = PP[2][10];
wire sF1i2L12, cF1i2L12;
FA F1i2L12( sF1i2L12,cF1i2L12,F1i2L12_inp1,F1i2L12_inp2,F1i2L12_inp3 );

wire F2i2L12_inp1, F2i2L12_inp2, F2i2L12_inp3;
assign F2i2L12_inp1 = PP[3][9];
assign F2i2L12_inp2 = PP[4][8];
assign F2i2L12_inp3 = PP[5][7];
wire sF2i2L12, cF2i2L12;
FA F2i2L12( sF2i2L12,cF2i2L12,F2i2L12_inp1,F2i2L12_inp2,F2i2L12_inp3 );

wire F3i2L12_inp1, F3i2L12_inp2, F3i2L12_inp3;
assign F3i2L12_inp1 = PP[6][6];
assign F3i2L12_inp2 = PP[7][5];
assign F3i2L12_inp3 = PP[8][4];
wire sF3i2L12, cF3i2L12;
FA F3i2L12( sF3i2L12,cF3i2L12,F3i2L12_inp1,F3i2L12_inp2,F3i2L12_inp3 );

wire Hi2L12_inp1, Hi2L12_inp2;
assign Hi2L12_inp1 = PP[9][3];
assign Hi2L12_inp2 = PP[10][2];
wire sHi2L12, cHi2L12;
HA Hi2L12 ( sHi2L12,cHi2L12,Hi2L12_inp1,Hi2L12_inp2 );

wire F1i2L13_inp1, F1i2L13_inp2, F1i2L13_inp3;
assign F1i2L13_inp1 = PP[3][10];
assign F1i2L13_inp2 = PP[4][9];
assign F1i2L13_inp3 = PP[5][8];
wire sF1i2L13, cF1i2L13;
FA F1i2L13( sF1i2L13,cF1i2L13,F1i2L13_inp1,F1i2L13_inp2,F1i2L13_inp3 );

wire F2i2L13_inp1, F2i2L13_inp2, F2i2L13_inp3;
assign F2i2L13_inp1 = PP[6][7];
assign F2i2L13_inp2 = PP[7][6];
assign F2i2L13_inp3 = PP[8][5];
wire sF2i2L13, cF2i2L13;
FA F2i2L13( sF2i2L13,cF2i2L13,F2i2L13_inp1,F2i2L13_inp2,F2i2L13_inp3 );

wire F3i2L13_inp1, F3i2L13_inp2, F3i2L13_inp3;
assign F3i2L13_inp1 = PP[9][4];
assign F3i2L13_inp2 = PP[10][3];
assign F3i2L13_inp3 = PP[11][2];
wire sF3i2L13, cF3i2L13;
FA F3i2L13( sF3i2L13,cF3i2L13,F3i2L13_inp1,F3i2L13_inp2,F3i2L13_inp3 );

wire F4i2L13_inp1, F4i2L13_inp2, F4i2L13_inp3;
assign F4i2L13_inp1 = PP[12][1];
assign F4i2L13_inp2 = PP[13][0];
assign F4i2L13_inp3 = CV[13];
wire sF4i2L13, cF4i2L13;
FA F4i2L13( sF4i2L13,cF4i2L13,F4i2L13_inp1,F4i2L13_inp2,F4i2L13_inp3 );

wire F1i2L14_inp1, F1i2L14_inp2, F1i2L14_inp3;
assign F1i2L14_inp1 = PP[4][10];
assign F1i2L14_inp2 = PP[5][9];
assign F1i2L14_inp3 = PP[6][8];
wire sF1i2L14, cF1i2L14;
FA F1i2L14( sF1i2L14,cF1i2L14,F1i2L14_inp1,F1i2L14_inp2,F1i2L14_inp3 );

wire F2i2L14_inp1, F2i2L14_inp2, F2i2L14_inp3;
assign F2i2L14_inp1 = PP[7][7];
assign F2i2L14_inp2 = PP[8][6];
assign F2i2L14_inp3 = PP[9][5];
wire sF2i2L14, cF2i2L14;
FA F2i2L14( sF2i2L14,cF2i2L14,F2i2L14_inp1,F2i2L14_inp2,F2i2L14_inp3 );

wire F3i2L14_inp1, F3i2L14_inp2, F3i2L14_inp3;
assign F3i2L14_inp1 = PP[10][4];
assign F3i2L14_inp2 = PP[11][3];
assign F3i2L14_inp3 = PP[12][2];
wire sF3i2L14, cF3i2L14;
FA F3i2L14( sF3i2L14,cF3i2L14,F3i2L14_inp1,F3i2L14_inp2,F3i2L14_inp3 );

wire F4i2L14_inp1, F4i2L14_inp2, F4i2L14_inp3;
assign F4i2L14_inp1 = PP[13][1];
assign F4i2L14_inp2 = PP[14][0];
assign F4i2L14_inp3 = cF1i1L13;
wire sF4i2L14, cF4i2L14;
FA F4i2L14( sF4i2L14,cF4i2L14,F4i2L14_inp1,F4i2L14_inp2,F4i2L14_inp3 );

wire F1i2L15_inp1, F1i2L15_inp2, F1i2L15_inp3;
assign F1i2L15_inp1 = PP[5][10];
assign F1i2L15_inp2 = PP[6][9];
assign F1i2L15_inp3 = PP[7][8];
wire sF1i2L15, cF1i2L15;
FA F1i2L15( sF1i2L15,cF1i2L15,F1i2L15_inp1,F1i2L15_inp2,F1i2L15_inp3 );

wire F2i2L15_inp1, F2i2L15_inp2, F2i2L15_inp3;
assign F2i2L15_inp1 = PP[8][7];
assign F2i2L15_inp2 = PP[9][6];
assign F2i2L15_inp3 = PP[10][5];
wire sF2i2L15, cF2i2L15;
FA F2i2L15( sF2i2L15,cF2i2L15,F2i2L15_inp1,F2i2L15_inp2,F2i2L15_inp3 );

wire F3i2L15_inp1, F3i2L15_inp2, F3i2L15_inp3;
assign F3i2L15_inp1 = PP[11][4];
assign F3i2L15_inp2 = PP[12][3];
assign F3i2L15_inp3 = PP[13][2];
wire sF3i2L15, cF3i2L15;
FA F3i2L15( sF3i2L15,cF3i2L15,F3i2L15_inp1,F3i2L15_inp2,F3i2L15_inp3 );

wire F4i2L15_inp1, F4i2L15_inp2, F4i2L15_inp3;
assign F4i2L15_inp1 = PP[14][1];
assign F4i2L15_inp2 = PP[15][0];
assign F4i2L15_inp3 = cF1i1L14;
wire sF4i2L15, cF4i2L15;
FA F4i2L15( sF4i2L15,cF4i2L15,F4i2L15_inp1,F4i2L15_inp2,F4i2L15_inp3 );

wire F1i2L16_inp1, F1i2L16_inp2, F1i2L16_inp3;
assign F1i2L16_inp1 = PP[5][11];
assign F1i2L16_inp2 = PP[6][10];
assign F1i2L16_inp3 = PP[7][9];
wire sF1i2L16, cF1i2L16;
FA F1i2L16( sF1i2L16,cF1i2L16,F1i2L16_inp1,F1i2L16_inp2,F1i2L16_inp3 );

wire F2i2L16_inp1, F2i2L16_inp2, F2i2L16_inp3;
assign F2i2L16_inp1 = PP[8][8];
assign F2i2L16_inp2 = PP[9][7];
assign F2i2L16_inp3 = PP[10][6];
wire sF2i2L16, cF2i2L16;
FA F2i2L16( sF2i2L16,cF2i2L16,F2i2L16_inp1,F2i2L16_inp2,F2i2L16_inp3 );

wire F3i2L16_inp1, F3i2L16_inp2, F3i2L16_inp3;
assign F3i2L16_inp1 = PP[11][5];
assign F3i2L16_inp2 = PP[12][4];
assign F3i2L16_inp3 = PP[13][3];
wire sF3i2L16, cF3i2L16;
FA F3i2L16( sF3i2L16,cF3i2L16,F3i2L16_inp1,F3i2L16_inp2,F3i2L16_inp3 );

wire F4i2L16_inp1, F4i2L16_inp2, F4i2L16_inp3;
assign F4i2L16_inp1 = PP[14][2];
assign F4i2L16_inp2 = PP[15][1];
assign F4i2L16_inp3 = cF1i1L15;
wire sF4i2L16, cF4i2L16;
FA F4i2L16( sF4i2L16,cF4i2L16,F4i2L16_inp1,F4i2L16_inp2,F4i2L16_inp3 );

wire F1i2L17_inp1, F1i2L17_inp2, F1i2L17_inp3;
assign F1i2L17_inp1 = ~PP[4][13];
assign F1i2L17_inp2 = PP[5][12];
assign F1i2L17_inp3 = PP[6][11];
wire sF1i2L17, cF1i2L17;
FA F1i2L17( sF1i2L17,cF1i2L17,F1i2L17_inp1,F1i2L17_inp2,F1i2L17_inp3 );

wire F2i2L17_inp1, F2i2L17_inp2, F2i2L17_inp3;
assign F2i2L17_inp1 = PP[7][10];
assign F2i2L17_inp2 = PP[8][9];
assign F2i2L17_inp3 = PP[9][8];
wire sF2i2L17, cF2i2L17;
FA F2i2L17( sF2i2L17,cF2i2L17,F2i2L17_inp1,F2i2L17_inp2,F2i2L17_inp3 );

wire F3i2L17_inp1, F3i2L17_inp2, F3i2L17_inp3;
assign F3i2L17_inp1 = PP[10][7];
assign F3i2L17_inp2 = PP[11][6];
assign F3i2L17_inp3 = PP[12][5];
wire sF3i2L17, cF3i2L17;
FA F3i2L17( sF3i2L17,cF3i2L17,F3i2L17_inp1,F3i2L17_inp2,F3i2L17_inp3 );

wire F4i2L17_inp1, F4i2L17_inp2, F4i2L17_inp3;
assign F4i2L17_inp1 = PP[13][4];
assign F4i2L17_inp2 = PP[14][3];
assign F4i2L17_inp3 = PP[15][2];
wire sF4i2L17, cF4i2L17;
FA F4i2L17( sF4i2L17,cF4i2L17,F4i2L17_inp1,F4i2L17_inp2,F4i2L17_inp3 );

wire F1i2L18_inp1, F1i2L18_inp2, F1i2L18_inp3;
assign F1i2L18_inp1 = ~PP[5][13];
assign F1i2L18_inp2 = PP[6][12];
assign F1i2L18_inp3 = PP[7][11];
wire sF1i2L18, cF1i2L18;
FA F1i2L18( sF1i2L18,cF1i2L18,F1i2L18_inp1,F1i2L18_inp2,F1i2L18_inp3 );

wire F2i2L18_inp1, F2i2L18_inp2, F2i2L18_inp3;
assign F2i2L18_inp1 = PP[8][10];
assign F2i2L18_inp2 = PP[9][9];
assign F2i2L18_inp3 = PP[10][8];
wire sF2i2L18, cF2i2L18;
FA F2i2L18( sF2i2L18,cF2i2L18,F2i2L18_inp1,F2i2L18_inp2,F2i2L18_inp3 );

wire F3i2L18_inp1, F3i2L18_inp2, F3i2L18_inp3;
assign F3i2L18_inp1 = PP[11][7];
assign F3i2L18_inp2 = PP[12][6];
assign F3i2L18_inp3 = PP[13][5];
wire sF3i2L18, cF3i2L18;
FA F3i2L18( sF3i2L18,cF3i2L18,F3i2L18_inp1,F3i2L18_inp2,F3i2L18_inp3 );

wire F1i2L19_inp1, F1i2L19_inp2, F1i2L19_inp3;
assign F1i2L19_inp1 = ~PP[6][13];
assign F1i2L19_inp2 = PP[7][12];
assign F1i2L19_inp3 = PP[8][11];
wire sF1i2L19, cF1i2L19;
FA F1i2L19( sF1i2L19,cF1i2L19,F1i2L19_inp1,F1i2L19_inp2,F1i2L19_inp3 );

wire F2i2L19_inp1, F2i2L19_inp2, F2i2L19_inp3;
assign F2i2L19_inp1 = PP[9][10];
assign F2i2L19_inp2 = PP[10][9];
assign F2i2L19_inp3 = PP[11][8];
wire sF2i2L19, cF2i2L19;
FA F2i2L19( sF2i2L19,cF2i2L19,F2i2L19_inp1,F2i2L19_inp2,F2i2L19_inp3 );

wire F1i2L20_inp1, F1i2L20_inp2, F1i2L20_inp3;
assign F1i2L20_inp1 = ~PP[7][13];
assign F1i2L20_inp2 = PP[8][12];
assign F1i2L20_inp3 = PP[9][11];
wire sF1i2L20, cF1i2L20;
FA F1i2L20( sF1i2L20,cF1i2L20,F1i2L20_inp1,F1i2L20_inp2,F1i2L20_inp3 );



///////////// Iteration Number =3///////////////////





wire Hi3L6_inp1, Hi3L6_inp2;
assign Hi3L6_inp1 = PP[0][6];
assign Hi3L6_inp2 = PP[1][5];
wire sHi3L6, cHi3L6;
HA Hi3L6 ( sHi3L6,cHi3L6,Hi3L6_inp1,Hi3L6_inp2 );

wire F1i3L7_inp1, F1i3L7_inp2, F1i3L7_inp3;
assign F1i3L7_inp1 = PP[0][7];
assign F1i3L7_inp2 = PP[1][6];
assign F1i3L7_inp3 = PP[2][5];
wire sF1i3L7, cF1i3L7;
FA F1i3L7( sF1i3L7,cF1i3L7,F1i3L7_inp1,F1i3L7_inp2,F1i3L7_inp3 );

wire Hi3L7_inp1, Hi3L7_inp2;
assign Hi3L7_inp1 = PP[3][4];
assign Hi3L7_inp2 = PP[4][3];
wire sHi3L7, cHi3L7;
HA Hi3L7 ( sHi3L7,cHi3L7,Hi3L7_inp1,Hi3L7_inp2 );

wire F1i3L8_inp1, F1i3L8_inp2, F1i3L8_inp3;
assign F1i3L8_inp1 = PP[0][8];
assign F1i3L8_inp2 = PP[1][7];
assign F1i3L8_inp3 = PP[2][6];
wire sF1i3L8, cF1i3L8;
FA F1i3L8( sF1i3L8,cF1i3L8,F1i3L8_inp1,F1i3L8_inp2,F1i3L8_inp3 );

wire F2i3L8_inp1, F2i3L8_inp2, F2i3L8_inp3;
assign F2i3L8_inp1 = PP[3][5];
assign F2i3L8_inp2 = PP[4][4];
assign F2i3L8_inp3 = PP[5][3];
wire sF2i3L8, cF2i3L8;
FA F2i3L8( sF2i3L8,cF2i3L8,F2i3L8_inp1,F2i3L8_inp2,F2i3L8_inp3 );

wire Hi3L8_inp1, Hi3L8_inp2;
assign Hi3L8_inp1 = PP[6][2];
assign Hi3L8_inp2 = PP[7][1];
wire sHi3L8, cHi3L8;
HA Hi3L8 ( sHi3L8,cHi3L8,Hi3L8_inp1,Hi3L8_inp2 );

wire F1i3L9_inp1, F1i3L9_inp2, F1i3L9_inp3;
assign F1i3L9_inp1 = PP[2][7];
assign F1i3L9_inp2 = PP[3][6];
assign F1i3L9_inp3 = PP[4][5];
wire sF1i3L9, cF1i3L9;
FA F1i3L9( sF1i3L9,cF1i3L9,F1i3L9_inp1,F1i3L9_inp2,F1i3L9_inp3 );

wire F2i3L9_inp1, F2i3L9_inp2, F2i3L9_inp3;
assign F2i3L9_inp1 = PP[5][4];
assign F2i3L9_inp2 = PP[6][3];
assign F2i3L9_inp3 = PP[7][2];
wire sF2i3L9, cF2i3L9;
FA F2i3L9( sF2i3L9,cF2i3L9,F2i3L9_inp1,F2i3L9_inp2,F2i3L9_inp3 );

wire F3i3L9_inp1, F3i3L9_inp2, F3i3L9_inp3;
assign F3i3L9_inp1 = PP[8][1];
assign F3i3L9_inp2 = PP[9][0];
assign F3i3L9_inp3 = sHi2L9;
wire sF3i3L9, cF3i3L9;
FA F3i3L9( sF3i3L9,cF3i3L9,F3i3L9_inp1,F3i3L9_inp2,F3i3L9_inp3 );

wire F1i3L10_inp1, F1i3L10_inp2, F1i3L10_inp3;
assign F1i3L10_inp1 = PP[5][5];
assign F1i3L10_inp2 = PP[6][4];
assign F1i3L10_inp3 = PP[7][3];
wire sF1i3L10, cF1i3L10;
FA F1i3L10( sF1i3L10,cF1i3L10,F1i3L10_inp1,F1i3L10_inp2,F1i3L10_inp3 );

wire F2i3L10_inp1, F2i3L10_inp2, F2i3L10_inp3;
assign F2i3L10_inp1 = PP[8][2];
assign F2i3L10_inp2 = PP[9][1];
assign F2i3L10_inp3 = PP[10][0];
wire sF2i3L10, cF2i3L10;
FA F2i3L10( sF2i3L10,cF2i3L10,F2i3L10_inp1,F2i3L10_inp2,F2i3L10_inp3 );

wire F3i3L10_inp1, F3i3L10_inp2, F3i3L10_inp3;
assign F3i3L10_inp1 = cHi2L9;
assign F3i3L10_inp2 = sF1i2L10;
assign F3i3L10_inp3 = sHi2L10;
wire sF3i3L10, cF3i3L10;
FA F3i3L10( sF3i3L10,cF3i3L10,F3i3L10_inp1,F3i3L10_inp2,F3i3L10_inp3 );

wire F1i3L11_inp1, F1i3L11_inp2, F1i3L11_inp3;
assign F1i3L11_inp1 = PP[8][3];
assign F1i3L11_inp2 = PP[9][2];
assign F1i3L11_inp3 = PP[10][1];
wire sF1i3L11, cF1i3L11;
FA F1i3L11( sF1i3L11,cF1i3L11,F1i3L11_inp1,F1i3L11_inp2,F1i3L11_inp3 );

wire F2i3L11_inp1, F2i3L11_inp2, F2i3L11_inp3;
assign F2i3L11_inp1 = PP[11][0];
assign F2i3L11_inp2 = cF1i2L10;
assign F2i3L11_inp3 = cHi2L10;
wire sF2i3L11, cF2i3L11;
FA F2i3L11( sF2i3L11,cF2i3L11,F2i3L11_inp1,F2i3L11_inp2,F2i3L11_inp3 );

wire F3i3L11_inp1, F3i3L11_inp2, F3i3L11_inp3;
assign F3i3L11_inp1 = sF1i2L11;
assign F3i3L11_inp2 = sF2i2L11;
assign F3i3L11_inp3 = sHi2L11;
wire sF3i3L11, cF3i3L11;
FA F3i3L11( sF3i3L11,cF3i3L11,F3i3L11_inp1,F3i3L11_inp2,F3i3L11_inp3 );

wire F1i3L12_inp1, F1i3L12_inp2, F1i3L12_inp3;
assign F1i3L12_inp1 = PP[11][1];
assign F1i3L12_inp2 = PP[12][0];
assign F1i3L12_inp3 = cF1i2L11;
wire sF1i3L12, cF1i3L12;
FA F1i3L12( sF1i3L12,cF1i3L12,F1i3L12_inp1,F1i3L12_inp2,F1i3L12_inp3 );

wire F2i3L12_inp1, F2i3L12_inp2, F2i3L12_inp3;
assign F2i3L12_inp1 = cF2i2L11;
assign F2i3L12_inp2 = cHi2L11;
assign F2i3L12_inp3 = sF1i2L12;
wire sF2i3L12, cF2i3L12;
FA F2i3L12( sF2i3L12,cF2i3L12,F2i3L12_inp1,F2i3L12_inp2,F2i3L12_inp3 );

wire F3i3L12_inp1, F3i3L12_inp2, F3i3L12_inp3;
assign F3i3L12_inp1 = sF2i2L12;
assign F3i3L12_inp2 = sF3i2L12;
assign F3i3L12_inp3 = sHi2L12;
wire sF3i3L12, cF3i3L12;
FA F3i3L12( sF3i3L12,cF3i3L12,F3i3L12_inp1,F3i3L12_inp2,F3i3L12_inp3 );

wire F1i3L13_inp1, F1i3L13_inp2, F1i3L13_inp3;
assign F1i3L13_inp1 = sF1i1L13;
assign F1i3L13_inp2 = cF1i2L12;
assign F1i3L13_inp3 = cF2i2L12;
wire sF1i3L13, cF1i3L13;
FA F1i3L13( sF1i3L13,cF1i3L13,F1i3L13_inp1,F1i3L13_inp2,F1i3L13_inp3 );

wire F2i3L13_inp1, F2i3L13_inp2, F2i3L13_inp3;
assign F2i3L13_inp1 = cF3i2L12;
assign F2i3L13_inp2 = cHi2L12;
assign F2i3L13_inp3 = sF1i2L13;
wire sF2i3L13, cF2i3L13;
FA F2i3L13( sF2i3L13,cF2i3L13,F2i3L13_inp1,F2i3L13_inp2,F2i3L13_inp3 );

wire F3i3L13_inp1, F3i3L13_inp2, F3i3L13_inp3;
assign F3i3L13_inp1 = sF2i2L13;
assign F3i3L13_inp2 = sF3i2L13;
assign F3i3L13_inp3 = sF4i2L13;
wire sF3i3L13, cF3i3L13;
FA F3i3L13( sF3i3L13,cF3i3L13,F3i3L13_inp1,F3i3L13_inp2,F3i3L13_inp3 );

wire F1i3L14_inp1, F1i3L14_inp2, F1i3L14_inp3;
assign F1i3L14_inp1 = sF1i1L14;
assign F1i3L14_inp2 = cF1i2L13;
assign F1i3L14_inp3 = cF2i2L13;
wire sF1i3L14, cF1i3L14;
FA F1i3L14( sF1i3L14,cF1i3L14,F1i3L14_inp1,F1i3L14_inp2,F1i3L14_inp3 );

wire F2i3L14_inp1, F2i3L14_inp2, F2i3L14_inp3;
assign F2i3L14_inp1 = cF3i2L13;
assign F2i3L14_inp2 = cF4i2L13;
assign F2i3L14_inp3 = sF1i2L14;
wire sF2i3L14, cF2i3L14;
FA F2i3L14( sF2i3L14,cF2i3L14,F2i3L14_inp1,F2i3L14_inp2,F2i3L14_inp3 );

wire F3i3L14_inp1, F3i3L14_inp2, F3i3L14_inp3;
assign F3i3L14_inp1 = sF2i2L14;
assign F3i3L14_inp2 = sF3i2L14;
assign F3i3L14_inp3 = sF4i2L14;
wire sF3i3L14, cF3i3L14;
FA F3i3L14( sF3i3L14,cF3i3L14,F3i3L14_inp1,F3i3L14_inp2,F3i3L14_inp3 );

wire F1i3L15_inp1, F1i3L15_inp2, F1i3L15_inp3;
assign F1i3L15_inp1 = sF1i1L15;
assign F1i3L15_inp2 = cF1i2L14;
assign F1i3L15_inp3 = cF2i2L14;
wire sF1i3L15, cF1i3L15;
FA F1i3L15( sF1i3L15,cF1i3L15,F1i3L15_inp1,F1i3L15_inp2,F1i3L15_inp3 );

wire F2i3L15_inp1, F2i3L15_inp2, F2i3L15_inp3;
assign F2i3L15_inp1 = cF3i2L14;
assign F2i3L15_inp2 = cF4i2L14;
assign F2i3L15_inp3 = sF1i2L15;
wire sF2i3L15, cF2i3L15;
FA F2i3L15( sF2i3L15,cF2i3L15,F2i3L15_inp1,F2i3L15_inp2,F2i3L15_inp3 );

wire F3i3L15_inp1, F3i3L15_inp2, F3i3L15_inp3;
assign F3i3L15_inp1 = sF2i2L15;
assign F3i3L15_inp2 = sF3i2L15;
assign F3i3L15_inp3 = sF4i2L15;
wire sF3i3L15, cF3i3L15;
FA F3i3L15( sF3i3L15,cF3i3L15,F3i3L15_inp1,F3i3L15_inp2,F3i3L15_inp3 );

wire F1i3L16_inp1, F1i3L16_inp2, F1i3L16_inp3;
assign F1i3L16_inp1 = sHi1L16;
assign F1i3L16_inp2 = cF1i2L15;
assign F1i3L16_inp3 = cF2i2L15;
wire sF1i3L16, cF1i3L16;
FA F1i3L16( sF1i3L16,cF1i3L16,F1i3L16_inp1,F1i3L16_inp2,F1i3L16_inp3 );

wire F2i3L16_inp1, F2i3L16_inp2, F2i3L16_inp3;
assign F2i3L16_inp1 = cF3i2L15;
assign F2i3L16_inp2 = cF4i2L15;
assign F2i3L16_inp3 = sF1i2L16;
wire sF2i3L16, cF2i3L16;
FA F2i3L16( sF2i3L16,cF2i3L16,F2i3L16_inp1,F2i3L16_inp2,F2i3L16_inp3 );

wire F3i3L16_inp1, F3i3L16_inp2, F3i3L16_inp3;
assign F3i3L16_inp1 = sF2i2L16;
assign F3i3L16_inp2 = sF3i2L16;
assign F3i3L16_inp3 = sF4i2L16;
wire sF3i3L16, cF3i3L16;
FA F3i3L16( sF3i3L16,cF3i3L16,F3i3L16_inp1,F3i3L16_inp2,F3i3L16_inp3 );

wire F1i3L17_inp1, F1i3L17_inp2, F1i3L17_inp3;
assign F1i3L17_inp1 = cHi1L16;
assign F1i3L17_inp2 = cF1i2L16;
assign F1i3L17_inp3 = cF2i2L16;
wire sF1i3L17, cF1i3L17;
FA F1i3L17( sF1i3L17,cF1i3L17,F1i3L17_inp1,F1i3L17_inp2,F1i3L17_inp3 );

wire F2i3L17_inp1, F2i3L17_inp2, F2i3L17_inp3;
assign F2i3L17_inp1 = cF3i2L16;
assign F2i3L17_inp2 = cF4i2L16;
assign F2i3L17_inp3 = sF1i2L17;
wire sF2i3L17, cF2i3L17;
FA F2i3L17( sF2i3L17,cF2i3L17,F2i3L17_inp1,F2i3L17_inp2,F2i3L17_inp3 );

wire F3i3L17_inp1, F3i3L17_inp2, F3i3L17_inp3;
assign F3i3L17_inp1 = sF2i2L17;
assign F3i3L17_inp2 = sF3i2L17;
assign F3i3L17_inp3 = sF4i2L17;
wire sF3i3L17, cF3i3L17;
FA F3i3L17( sF3i3L17,cF3i3L17,F3i3L17_inp1,F3i3L17_inp2,F3i3L17_inp3 );

wire F1i3L18_inp1, F1i3L18_inp2, F1i3L18_inp3;
assign F1i3L18_inp1 = PP[14][4];
assign F1i3L18_inp2 = PP[15][3];
assign F1i3L18_inp3 = cF1i2L17;
wire sF1i3L18, cF1i3L18;
FA F1i3L18( sF1i3L18,cF1i3L18,F1i3L18_inp1,F1i3L18_inp2,F1i3L18_inp3 );

wire F2i3L18_inp1, F2i3L18_inp2, F2i3L18_inp3;
assign F2i3L18_inp1 = cF2i2L17;
assign F2i3L18_inp2 = cF3i2L17;
assign F2i3L18_inp3 = cF4i2L17;
wire sF2i3L18, cF2i3L18;
FA F2i3L18( sF2i3L18,cF2i3L18,F2i3L18_inp1,F2i3L18_inp2,F2i3L18_inp3 );

wire F3i3L18_inp1, F3i3L18_inp2, F3i3L18_inp3;
assign F3i3L18_inp1 = sF1i2L18;
assign F3i3L18_inp2 = sF2i2L18;
assign F3i3L18_inp3 = sF3i2L18;
wire sF3i3L18, cF3i3L18;
FA F3i3L18( sF3i3L18,cF3i3L18,F3i3L18_inp1,F3i3L18_inp2,F3i3L18_inp3 );

wire F1i3L19_inp1, F1i3L19_inp2, F1i3L19_inp3;
assign F1i3L19_inp1 = PP[12][7];
assign F1i3L19_inp2 = PP[13][6];
assign F1i3L19_inp3 = PP[14][5];
wire sF1i3L19, cF1i3L19;
FA F1i3L19( sF1i3L19,cF1i3L19,F1i3L19_inp1,F1i3L19_inp2,F1i3L19_inp3 );

wire F2i3L19_inp1, F2i3L19_inp2, F2i3L19_inp3;
assign F2i3L19_inp1 = PP[15][4];
assign F2i3L19_inp2 = cF1i2L18;
assign F2i3L19_inp3 = cF2i2L18;
wire sF2i3L19, cF2i3L19;
FA F2i3L19( sF2i3L19,cF2i3L19,F2i3L19_inp1,F2i3L19_inp2,F2i3L19_inp3 );

wire F3i3L19_inp1, F3i3L19_inp2, F3i3L19_inp3;
assign F3i3L19_inp1 = cF3i2L18;
assign F3i3L19_inp2 = sF1i2L19;
assign F3i3L19_inp3 = sF2i2L19;
wire sF3i3L19, cF3i3L19;
FA F3i3L19( sF3i3L19,cF3i3L19,F3i3L19_inp1,F3i3L19_inp2,F3i3L19_inp3 );

wire F1i3L20_inp1, F1i3L20_inp2, F1i3L20_inp3;
assign F1i3L20_inp1 = PP[10][10];
assign F1i3L20_inp2 = PP[11][9];
assign F1i3L20_inp3 = PP[12][8];
wire sF1i3L20, cF1i3L20;
FA F1i3L20( sF1i3L20,cF1i3L20,F1i3L20_inp1,F1i3L20_inp2,F1i3L20_inp3 );

wire F2i3L20_inp1, F2i3L20_inp2, F2i3L20_inp3;
assign F2i3L20_inp1 = PP[13][7];
assign F2i3L20_inp2 = PP[14][6];
assign F2i3L20_inp3 = PP[15][5];
wire sF2i3L20, cF2i3L20;
FA F2i3L20( sF2i3L20,cF2i3L20,F2i3L20_inp1,F2i3L20_inp2,F2i3L20_inp3 );

wire F3i3L20_inp1, F3i3L20_inp2, F3i3L20_inp3;
assign F3i3L20_inp1 = cF1i2L19;
assign F3i3L20_inp2 = cF2i2L19;
assign F3i3L20_inp3 = sF1i2L20;
wire sF3i3L20, cF3i3L20;
FA F3i3L20( sF3i3L20,cF3i3L20,F3i3L20_inp1,F3i3L20_inp2,F3i3L20_inp3 );

wire F1i3L21_inp1, F1i3L21_inp2, F1i3L21_inp3;
assign F1i3L21_inp1 = ~PP[8][13];
assign F1i3L21_inp2 = PP[9][12];
assign F1i3L21_inp3 = PP[10][11];
wire sF1i3L21, cF1i3L21;
FA F1i3L21( sF1i3L21,cF1i3L21,F1i3L21_inp1,F1i3L21_inp2,F1i3L21_inp3 );

wire F2i3L21_inp1, F2i3L21_inp2, F2i3L21_inp3;
assign F2i3L21_inp1 = PP[11][10];
assign F2i3L21_inp2 = PP[12][9];
assign F2i3L21_inp3 = PP[13][8];
wire sF2i3L21, cF2i3L21;
FA F2i3L21( sF2i3L21,cF2i3L21,F2i3L21_inp1,F2i3L21_inp2,F2i3L21_inp3 );

wire F3i3L21_inp1, F3i3L21_inp2, F3i3L21_inp3;
assign F3i3L21_inp1 = PP[14][7];
assign F3i3L21_inp2 = PP[15][6];
assign F3i3L21_inp3 = cF1i2L20;
wire sF3i3L21, cF3i3L21;
FA F3i3L21( sF3i3L21,cF3i3L21,F3i3L21_inp1,F3i3L21_inp2,F3i3L21_inp3 );

wire F1i3L22_inp1, F1i3L22_inp2, F1i3L22_inp3;
assign F1i3L22_inp1 = ~PP[9][13];
assign F1i3L22_inp2 = PP[10][12];
assign F1i3L22_inp3 = PP[11][11];
wire sF1i3L22, cF1i3L22;
FA F1i3L22( sF1i3L22,cF1i3L22,F1i3L22_inp1,F1i3L22_inp2,F1i3L22_inp3 );

wire F2i3L22_inp1, F2i3L22_inp2, F2i3L22_inp3;
assign F2i3L22_inp1 = PP[12][10];
assign F2i3L22_inp2 = PP[13][9];
assign F2i3L22_inp3 = PP[14][8];
wire sF2i3L22, cF2i3L22;
FA F2i3L22( sF2i3L22,cF2i3L22,F2i3L22_inp1,F2i3L22_inp2,F2i3L22_inp3 );

wire F1i3L23_inp1, F1i3L23_inp2, F1i3L23_inp3;
assign F1i3L23_inp1 = ~PP[10][13];
assign F1i3L23_inp2 = PP[11][12];
assign F1i3L23_inp3 = PP[12][11];
wire sF1i3L23, cF1i3L23;
FA F1i3L23( sF1i3L23,cF1i3L23,F1i3L23_inp1,F1i3L23_inp2,F1i3L23_inp3 );



///////////// Iteration Number =4///////////////////





wire Hi4L4_inp1, Hi4L4_inp2;
assign Hi4L4_inp1 = PP[0][4];
assign Hi4L4_inp2 = PP[1][3];
wire sHi4L4, cHi4L4;
HA Hi4L4 ( sHi4L4,cHi4L4,Hi4L4_inp1,Hi4L4_inp2 );

wire F1i4L5_inp1, F1i4L5_inp2, F1i4L5_inp3;
assign F1i4L5_inp1 = PP[0][5];
assign F1i4L5_inp2 = PP[1][4];
assign F1i4L5_inp3 = PP[2][3];
wire sF1i4L5, cF1i4L5;
FA F1i4L5( sF1i4L5,cF1i4L5,F1i4L5_inp1,F1i4L5_inp2,F1i4L5_inp3 );

wire Hi4L5_inp1, Hi4L5_inp2;
assign Hi4L5_inp1 = PP[3][2];
assign Hi4L5_inp2 = PP[4][1];
wire sHi4L5, cHi4L5;
HA Hi4L5 ( sHi4L5,cHi4L5,Hi4L5_inp1,Hi4L5_inp2 );

wire F1i4L6_inp1, F1i4L6_inp2, F1i4L6_inp3;
assign F1i4L6_inp1 = PP[2][4];
assign F1i4L6_inp2 = PP[3][3];
assign F1i4L6_inp3 = PP[4][2];
wire sF1i4L6, cF1i4L6;
FA F1i4L6( sF1i4L6,cF1i4L6,F1i4L6_inp1,F1i4L6_inp2,F1i4L6_inp3 );

wire F2i4L6_inp1, F2i4L6_inp2, F2i4L6_inp3;
assign F2i4L6_inp1 = PP[5][1];
assign F2i4L6_inp2 = PP[6][0];
assign F2i4L6_inp3 = sHi3L6;
wire sF2i4L6, cF2i4L6;
FA F2i4L6( sF2i4L6,cF2i4L6,F2i4L6_inp1,F2i4L6_inp2,F2i4L6_inp3 );

wire F1i4L7_inp1, F1i4L7_inp2, F1i4L7_inp3;
assign F1i4L7_inp1 = PP[5][2];
assign F1i4L7_inp2 = PP[6][1];
assign F1i4L7_inp3 = PP[7][0];
wire sF1i4L7, cF1i4L7;
FA F1i4L7( sF1i4L7,cF1i4L7,F1i4L7_inp1,F1i4L7_inp2,F1i4L7_inp3 );

wire F2i4L7_inp1, F2i4L7_inp2, F2i4L7_inp3;
assign F2i4L7_inp1 = cHi3L6;
assign F2i4L7_inp2 = sF1i3L7;
assign F2i4L7_inp3 = sHi3L7;
wire sF2i4L7, cF2i4L7;
FA F2i4L7( sF2i4L7,cF2i4L7,F2i4L7_inp1,F2i4L7_inp2,F2i4L7_inp3 );

wire F1i4L8_inp1, F1i4L8_inp2, F1i4L8_inp3;
assign F1i4L8_inp1 = PP[8][0];
assign F1i4L8_inp2 = cF1i3L7;
assign F1i4L8_inp3 = cHi3L7;
wire sF1i4L8, cF1i4L8;
FA F1i4L8( sF1i4L8,cF1i4L8,F1i4L8_inp1,F1i4L8_inp2,F1i4L8_inp3 );

wire F2i4L8_inp1, F2i4L8_inp2, F2i4L8_inp3;
assign F2i4L8_inp1 = sF1i3L8;
assign F2i4L8_inp2 = sF2i3L8;
assign F2i4L8_inp3 = sHi3L8;
wire sF2i4L8, cF2i4L8;
FA F2i4L8( sF2i4L8,cF2i4L8,F2i4L8_inp1,F2i4L8_inp2,F2i4L8_inp3 );

wire F1i4L9_inp1, F1i4L9_inp2, F1i4L9_inp3;
assign F1i4L9_inp1 = cF1i3L8;
assign F1i4L9_inp2 = cF2i3L8;
assign F1i4L9_inp3 = cHi3L8;
wire sF1i4L9, cF1i4L9;
FA F1i4L9( sF1i4L9,cF1i4L9,F1i4L9_inp1,F1i4L9_inp2,F1i4L9_inp3 );

wire F2i4L9_inp1, F2i4L9_inp2, F2i4L9_inp3;
assign F2i4L9_inp1 = sF1i3L9;
assign F2i4L9_inp2 = sF2i3L9;
assign F2i4L9_inp3 = sF3i3L9;
wire sF2i4L9, cF2i4L9;
FA F2i4L9( sF2i4L9,cF2i4L9,F2i4L9_inp1,F2i4L9_inp2,F2i4L9_inp3 );

wire F1i4L10_inp1, F1i4L10_inp2, F1i4L10_inp3;
assign F1i4L10_inp1 = cF1i3L9;
assign F1i4L10_inp2 = cF2i3L9;
assign F1i4L10_inp3 = cF3i3L9;
wire sF1i4L10, cF1i4L10;
FA F1i4L10( sF1i4L10,cF1i4L10,F1i4L10_inp1,F1i4L10_inp2,F1i4L10_inp3 );

wire F2i4L10_inp1, F2i4L10_inp2, F2i4L10_inp3;
assign F2i4L10_inp1 = sF1i3L10;
assign F2i4L10_inp2 = sF2i3L10;
assign F2i4L10_inp3 = sF3i3L10;
wire sF2i4L10, cF2i4L10;
FA F2i4L10( sF2i4L10,cF2i4L10,F2i4L10_inp1,F2i4L10_inp2,F2i4L10_inp3 );

wire F1i4L11_inp1, F1i4L11_inp2, F1i4L11_inp3;
assign F1i4L11_inp1 = cF1i3L10;
assign F1i4L11_inp2 = cF2i3L10;
assign F1i4L11_inp3 = cF3i3L10;
wire sF1i4L11, cF1i4L11;
FA F1i4L11( sF1i4L11,cF1i4L11,F1i4L11_inp1,F1i4L11_inp2,F1i4L11_inp3 );

wire F2i4L11_inp1, F2i4L11_inp2, F2i4L11_inp3;
assign F2i4L11_inp1 = sF1i3L11;
assign F2i4L11_inp2 = sF2i3L11;
assign F2i4L11_inp3 = sF3i3L11;
wire sF2i4L11, cF2i4L11;
FA F2i4L11( sF2i4L11,cF2i4L11,F2i4L11_inp1,F2i4L11_inp2,F2i4L11_inp3 );

wire F1i4L12_inp1, F1i4L12_inp2, F1i4L12_inp3;
assign F1i4L12_inp1 = cF1i3L11;
assign F1i4L12_inp2 = cF2i3L11;
assign F1i4L12_inp3 = cF3i3L11;
wire sF1i4L12, cF1i4L12;
FA F1i4L12( sF1i4L12,cF1i4L12,F1i4L12_inp1,F1i4L12_inp2,F1i4L12_inp3 );

wire F2i4L12_inp1, F2i4L12_inp2, F2i4L12_inp3;
assign F2i4L12_inp1 = sF1i3L12;
assign F2i4L12_inp2 = sF2i3L12;
assign F2i4L12_inp3 = sF3i3L12;
wire sF2i4L12, cF2i4L12;
FA F2i4L12( sF2i4L12,cF2i4L12,F2i4L12_inp1,F2i4L12_inp2,F2i4L12_inp3 );

wire F1i4L13_inp1, F1i4L13_inp2, F1i4L13_inp3;
assign F1i4L13_inp1 = cF1i3L12;
assign F1i4L13_inp2 = cF2i3L12;
assign F1i4L13_inp3 = cF3i3L12;
wire sF1i4L13, cF1i4L13;
FA F1i4L13( sF1i4L13,cF1i4L13,F1i4L13_inp1,F1i4L13_inp2,F1i4L13_inp3 );

wire F2i4L13_inp1, F2i4L13_inp2, F2i4L13_inp3;
assign F2i4L13_inp1 = sF1i3L13;
assign F2i4L13_inp2 = sF2i3L13;
assign F2i4L13_inp3 = sF3i3L13;
wire sF2i4L13, cF2i4L13;
FA F2i4L13( sF2i4L13,cF2i4L13,F2i4L13_inp1,F2i4L13_inp2,F2i4L13_inp3 );

wire F1i4L14_inp1, F1i4L14_inp2, F1i4L14_inp3;
assign F1i4L14_inp1 = cF1i3L13;
assign F1i4L14_inp2 = cF2i3L13;
assign F1i4L14_inp3 = cF3i3L13;
wire sF1i4L14, cF1i4L14;
FA F1i4L14( sF1i4L14,cF1i4L14,F1i4L14_inp1,F1i4L14_inp2,F1i4L14_inp3 );

wire F2i4L14_inp1, F2i4L14_inp2, F2i4L14_inp3;
assign F2i4L14_inp1 = sF1i3L14;
assign F2i4L14_inp2 = sF2i3L14;
assign F2i4L14_inp3 = sF3i3L14;
wire sF2i4L14, cF2i4L14;
FA F2i4L14( sF2i4L14,cF2i4L14,F2i4L14_inp1,F2i4L14_inp2,F2i4L14_inp3 );

wire F1i4L15_inp1, F1i4L15_inp2, F1i4L15_inp3;
assign F1i4L15_inp1 = cF1i3L14;
assign F1i4L15_inp2 = cF2i3L14;
assign F1i4L15_inp3 = cF3i3L14;
wire sF1i4L15, cF1i4L15;
FA F1i4L15( sF1i4L15,cF1i4L15,F1i4L15_inp1,F1i4L15_inp2,F1i4L15_inp3 );

wire F2i4L15_inp1, F2i4L15_inp2, F2i4L15_inp3;
assign F2i4L15_inp1 = sF1i3L15;
assign F2i4L15_inp2 = sF2i3L15;
assign F2i4L15_inp3 = sF3i3L15;
wire sF2i4L15, cF2i4L15;
FA F2i4L15( sF2i4L15,cF2i4L15,F2i4L15_inp1,F2i4L15_inp2,F2i4L15_inp3 );

wire F1i4L16_inp1, F1i4L16_inp2, F1i4L16_inp3;
assign F1i4L16_inp1 = cF1i3L15;
assign F1i4L16_inp2 = cF2i3L15;
assign F1i4L16_inp3 = cF3i3L15;
wire sF1i4L16, cF1i4L16;
FA F1i4L16( sF1i4L16,cF1i4L16,F1i4L16_inp1,F1i4L16_inp2,F1i4L16_inp3 );

wire F2i4L16_inp1, F2i4L16_inp2, F2i4L16_inp3;
assign F2i4L16_inp1 = sF1i3L16;
assign F2i4L16_inp2 = sF2i3L16;
assign F2i4L16_inp3 = sF3i3L16;
wire sF2i4L16, cF2i4L16;
FA F2i4L16( sF2i4L16,cF2i4L16,F2i4L16_inp1,F2i4L16_inp2,F2i4L16_inp3 );

wire F1i4L17_inp1, F1i4L17_inp2, F1i4L17_inp3;
assign F1i4L17_inp1 = cF1i3L16;
assign F1i4L17_inp2 = cF2i3L16;
assign F1i4L17_inp3 = cF3i3L16;
wire sF1i4L17, cF1i4L17;
FA F1i4L17( sF1i4L17,cF1i4L17,F1i4L17_inp1,F1i4L17_inp2,F1i4L17_inp3 );

wire F2i4L17_inp1, F2i4L17_inp2, F2i4L17_inp3;
assign F2i4L17_inp1 = sF1i3L17;
assign F2i4L17_inp2 = sF2i3L17;
assign F2i4L17_inp3 = sF3i3L17;
wire sF2i4L17, cF2i4L17;
FA F2i4L17( sF2i4L17,cF2i4L17,F2i4L17_inp1,F2i4L17_inp2,F2i4L17_inp3 );

wire F1i4L18_inp1, F1i4L18_inp2, F1i4L18_inp3;
assign F1i4L18_inp1 = cF1i3L17;
assign F1i4L18_inp2 = cF2i3L17;
assign F1i4L18_inp3 = cF3i3L17;
wire sF1i4L18, cF1i4L18;
FA F1i4L18( sF1i4L18,cF1i4L18,F1i4L18_inp1,F1i4L18_inp2,F1i4L18_inp3 );

wire F2i4L18_inp1, F2i4L18_inp2, F2i4L18_inp3;
assign F2i4L18_inp1 = sF1i3L18;
assign F2i4L18_inp2 = sF2i3L18;
assign F2i4L18_inp3 = sF3i3L18;
wire sF2i4L18, cF2i4L18;
FA F2i4L18( sF2i4L18,cF2i4L18,F2i4L18_inp1,F2i4L18_inp2,F2i4L18_inp3 );

wire F1i4L19_inp1, F1i4L19_inp2, F1i4L19_inp3;
assign F1i4L19_inp1 = cF1i3L18;
assign F1i4L19_inp2 = cF2i3L18;
assign F1i4L19_inp3 = cF3i3L18;
wire sF1i4L19, cF1i4L19;
FA F1i4L19( sF1i4L19,cF1i4L19,F1i4L19_inp1,F1i4L19_inp2,F1i4L19_inp3 );

wire F2i4L19_inp1, F2i4L19_inp2, F2i4L19_inp3;
assign F2i4L19_inp1 = sF1i3L19;
assign F2i4L19_inp2 = sF2i3L19;
assign F2i4L19_inp3 = sF3i3L19;
wire sF2i4L19, cF2i4L19;
FA F2i4L19( sF2i4L19,cF2i4L19,F2i4L19_inp1,F2i4L19_inp2,F2i4L19_inp3 );

wire F1i4L20_inp1, F1i4L20_inp2, F1i4L20_inp3;
assign F1i4L20_inp1 = cF1i3L19;
assign F1i4L20_inp2 = cF2i3L19;
assign F1i4L20_inp3 = cF3i3L19;
wire sF1i4L20, cF1i4L20;
FA F1i4L20( sF1i4L20,cF1i4L20,F1i4L20_inp1,F1i4L20_inp2,F1i4L20_inp3 );

wire F2i4L20_inp1, F2i4L20_inp2, F2i4L20_inp3;
assign F2i4L20_inp1 = sF1i3L20;
assign F2i4L20_inp2 = sF2i3L20;
assign F2i4L20_inp3 = sF3i3L20;
wire sF2i4L20, cF2i4L20;
FA F2i4L20( sF2i4L20,cF2i4L20,F2i4L20_inp1,F2i4L20_inp2,F2i4L20_inp3 );

wire F1i4L21_inp1, F1i4L21_inp2, F1i4L21_inp3;
assign F1i4L21_inp1 = cF1i3L20;
assign F1i4L21_inp2 = cF2i3L20;
assign F1i4L21_inp3 = cF3i3L20;
wire sF1i4L21, cF1i4L21;
FA F1i4L21( sF1i4L21,cF1i4L21,F1i4L21_inp1,F1i4L21_inp2,F1i4L21_inp3 );

wire F2i4L21_inp1, F2i4L21_inp2, F2i4L21_inp3;
assign F2i4L21_inp1 = sF1i3L21;
assign F2i4L21_inp2 = sF2i3L21;
assign F2i4L21_inp3 = sF3i3L21;
wire sF2i4L21, cF2i4L21;
FA F2i4L21( sF2i4L21,cF2i4L21,F2i4L21_inp1,F2i4L21_inp2,F2i4L21_inp3 );

wire F1i4L22_inp1, F1i4L22_inp2, F1i4L22_inp3;
assign F1i4L22_inp1 = PP[15][7];
assign F1i4L22_inp2 = cF1i3L21;
assign F1i4L22_inp3 = cF2i3L21;
wire sF1i4L22, cF1i4L22;
FA F1i4L22( sF1i4L22,cF1i4L22,F1i4L22_inp1,F1i4L22_inp2,F1i4L22_inp3 );

wire F2i4L22_inp1, F2i4L22_inp2, F2i4L22_inp3;
assign F2i4L22_inp1 = cF3i3L21;
assign F2i4L22_inp2 = sF1i3L22;
assign F2i4L22_inp3 = sF2i3L22;
wire sF2i4L22, cF2i4L22;
FA F2i4L22( sF2i4L22,cF2i4L22,F2i4L22_inp1,F2i4L22_inp2,F2i4L22_inp3 );

wire F1i4L23_inp1, F1i4L23_inp2, F1i4L23_inp3;
assign F1i4L23_inp1 = PP[13][10];
assign F1i4L23_inp2 = PP[14][9];
assign F1i4L23_inp3 = PP[15][8];
wire sF1i4L23, cF1i4L23;
FA F1i4L23( sF1i4L23,cF1i4L23,F1i4L23_inp1,F1i4L23_inp2,F1i4L23_inp3 );

wire F2i4L23_inp1, F2i4L23_inp2, F2i4L23_inp3;
assign F2i4L23_inp1 = cF1i3L22;
assign F2i4L23_inp2 = cF2i3L22;
assign F2i4L23_inp3 = sF1i3L23;
wire sF2i4L23, cF2i4L23;
FA F2i4L23( sF2i4L23,cF2i4L23,F2i4L23_inp1,F2i4L23_inp2,F2i4L23_inp3 );

wire F1i4L24_inp1, F1i4L24_inp2, F1i4L24_inp3;
assign F1i4L24_inp1 = ~PP[11][13];
assign F1i4L24_inp2 = PP[12][12];
assign F1i4L24_inp3 = PP[13][11];
wire sF1i4L24, cF1i4L24;
FA F1i4L24( sF1i4L24,cF1i4L24,F1i4L24_inp1,F1i4L24_inp2,F1i4L24_inp3 );

wire F2i4L24_inp1, F2i4L24_inp2, F2i4L24_inp3;
assign F2i4L24_inp1 = PP[14][10];
assign F2i4L24_inp2 = PP[15][9];
assign F2i4L24_inp3 = cF1i3L23;
wire sF2i4L24, cF2i4L24;
FA F2i4L24( sF2i4L24,cF2i4L24,F2i4L24_inp1,F2i4L24_inp2,F2i4L24_inp3 );

wire F1i4L25_inp1, F1i4L25_inp2, F1i4L25_inp3;
assign F1i4L25_inp1 = ~PP[12][13];
assign F1i4L25_inp2 = PP[13][12];
assign F1i4L25_inp3 = PP[14][11];
wire sF1i4L25, cF1i4L25;
FA F1i4L25( sF1i4L25,cF1i4L25,F1i4L25_inp1,F1i4L25_inp2,F1i4L25_inp3 );



///////////// Iteration Number =5///////////////////





wire Hi5L3_inp1, Hi5L3_inp2;
assign Hi5L3_inp1 = PP[0][3];
assign Hi5L3_inp2 = PP[1][2];
wire sHi5L3, cHi5L3;
HA Hi5L3 ( sHi5L3,cHi5L3,Hi5L3_inp1,Hi5L3_inp2 );

wire F1i5L4_inp1, F1i5L4_inp2, F1i5L4_inp3;
assign F1i5L4_inp1 = PP[2][2];
assign F1i5L4_inp2 = PP[3][1];
assign F1i5L4_inp3 = PP[4][0];
wire sF1i5L4, cF1i5L4;
FA F1i5L4( sF1i5L4,cF1i5L4,F1i5L4_inp1,F1i5L4_inp2,F1i5L4_inp3 );

wire F1i5L5_inp1, F1i5L5_inp2, F1i5L5_inp3;
assign F1i5L5_inp1 = PP[5][0];
assign F1i5L5_inp2 = cHi4L4;
assign F1i5L5_inp3 = sF1i4L5;
wire sF1i5L5, cF1i5L5;
FA F1i5L5( sF1i5L5,cF1i5L5,F1i5L5_inp1,F1i5L5_inp2,F1i5L5_inp3 );

wire F1i5L6_inp1, F1i5L6_inp2, F1i5L6_inp3;
assign F1i5L6_inp1 = cF1i4L5;
assign F1i5L6_inp2 = cHi4L5;
assign F1i5L6_inp3 = sF1i4L6;
wire sF1i5L6, cF1i5L6;
FA F1i5L6( sF1i5L6,cF1i5L6,F1i5L6_inp1,F1i5L6_inp2,F1i5L6_inp3 );

wire F1i5L7_inp1, F1i5L7_inp2, F1i5L7_inp3;
assign F1i5L7_inp1 = cF1i4L6;
assign F1i5L7_inp2 = cF2i4L6;
assign F1i5L7_inp3 = sF1i4L7;
wire sF1i5L7, cF1i5L7;
FA F1i5L7( sF1i5L7,cF1i5L7,F1i5L7_inp1,F1i5L7_inp2,F1i5L7_inp3 );

wire F1i5L8_inp1, F1i5L8_inp2, F1i5L8_inp3;
assign F1i5L8_inp1 = cF1i4L7;
assign F1i5L8_inp2 = cF2i4L7;
assign F1i5L8_inp3 = sF1i4L8;
wire sF1i5L8, cF1i5L8;
FA F1i5L8( sF1i5L8,cF1i5L8,F1i5L8_inp1,F1i5L8_inp2,F1i5L8_inp3 );

wire F1i5L9_inp1, F1i5L9_inp2, F1i5L9_inp3;
assign F1i5L9_inp1 = cF1i4L8;
assign F1i5L9_inp2 = cF2i4L8;
assign F1i5L9_inp3 = sF1i4L9;
wire sF1i5L9, cF1i5L9;
FA F1i5L9( sF1i5L9,cF1i5L9,F1i5L9_inp1,F1i5L9_inp2,F1i5L9_inp3 );

wire F1i5L10_inp1, F1i5L10_inp2, F1i5L10_inp3;
assign F1i5L10_inp1 = cF1i4L9;
assign F1i5L10_inp2 = cF2i4L9;
assign F1i5L10_inp3 = sF1i4L10;
wire sF1i5L10, cF1i5L10;
FA F1i5L10( sF1i5L10,cF1i5L10,F1i5L10_inp1,F1i5L10_inp2,F1i5L10_inp3 );

wire F1i5L11_inp1, F1i5L11_inp2, F1i5L11_inp3;
assign F1i5L11_inp1 = cF1i4L10;
assign F1i5L11_inp2 = cF2i4L10;
assign F1i5L11_inp3 = sF1i4L11;
wire sF1i5L11, cF1i5L11;
FA F1i5L11( sF1i5L11,cF1i5L11,F1i5L11_inp1,F1i5L11_inp2,F1i5L11_inp3 );

wire F1i5L12_inp1, F1i5L12_inp2, F1i5L12_inp3;
assign F1i5L12_inp1 = cF1i4L11;
assign F1i5L12_inp2 = cF2i4L11;
assign F1i5L12_inp3 = sF1i4L12;
wire sF1i5L12, cF1i5L12;
FA F1i5L12( sF1i5L12,cF1i5L12,F1i5L12_inp1,F1i5L12_inp2,F1i5L12_inp3 );

wire F1i5L13_inp1, F1i5L13_inp2, F1i5L13_inp3;
assign F1i5L13_inp1 = cF1i4L12;
assign F1i5L13_inp2 = cF2i4L12;
assign F1i5L13_inp3 = sF1i4L13;
wire sF1i5L13, cF1i5L13;
FA F1i5L13( sF1i5L13,cF1i5L13,F1i5L13_inp1,F1i5L13_inp2,F1i5L13_inp3 );

wire F1i5L14_inp1, F1i5L14_inp2, F1i5L14_inp3;
assign F1i5L14_inp1 = cF1i4L13;
assign F1i5L14_inp2 = cF2i4L13;
assign F1i5L14_inp3 = sF1i4L14;
wire sF1i5L14, cF1i5L14;
FA F1i5L14( sF1i5L14,cF1i5L14,F1i5L14_inp1,F1i5L14_inp2,F1i5L14_inp3 );

wire F1i5L15_inp1, F1i5L15_inp2, F1i5L15_inp3;
assign F1i5L15_inp1 = cF1i4L14;
assign F1i5L15_inp2 = cF2i4L14;
assign F1i5L15_inp3 = sF1i4L15;
wire sF1i5L15, cF1i5L15;
FA F1i5L15( sF1i5L15,cF1i5L15,F1i5L15_inp1,F1i5L15_inp2,F1i5L15_inp3 );

wire F1i5L16_inp1, F1i5L16_inp2, F1i5L16_inp3;
assign F1i5L16_inp1 = cF1i4L15;
assign F1i5L16_inp2 = cF2i4L15;
assign F1i5L16_inp3 = sF1i4L16;
wire sF1i5L16, cF1i5L16;
FA F1i5L16( sF1i5L16,cF1i5L16,F1i5L16_inp1,F1i5L16_inp2,F1i5L16_inp3 );

wire F1i5L17_inp1, F1i5L17_inp2, F1i5L17_inp3;
assign F1i5L17_inp1 = cF1i4L16;
assign F1i5L17_inp2 = cF2i4L16;
assign F1i5L17_inp3 = sF1i4L17;
wire sF1i5L17, cF1i5L17;
FA F1i5L17( sF1i5L17,cF1i5L17,F1i5L17_inp1,F1i5L17_inp2,F1i5L17_inp3 );

wire F1i5L18_inp1, F1i5L18_inp2, F1i5L18_inp3;
assign F1i5L18_inp1 = cF1i4L17;
assign F1i5L18_inp2 = cF2i4L17;
assign F1i5L18_inp3 = sF1i4L18;
wire sF1i5L18, cF1i5L18;
FA F1i5L18( sF1i5L18,cF1i5L18,F1i5L18_inp1,F1i5L18_inp2,F1i5L18_inp3 );

wire F1i5L19_inp1, F1i5L19_inp2, F1i5L19_inp3;
assign F1i5L19_inp1 = cF1i4L18;
assign F1i5L19_inp2 = cF2i4L18;
assign F1i5L19_inp3 = sF1i4L19;
wire sF1i5L19, cF1i5L19;
FA F1i5L19( sF1i5L19,cF1i5L19,F1i5L19_inp1,F1i5L19_inp2,F1i5L19_inp3 );

wire F1i5L20_inp1, F1i5L20_inp2, F1i5L20_inp3;
assign F1i5L20_inp1 = cF1i4L19;
assign F1i5L20_inp2 = cF2i4L19;
assign F1i5L20_inp3 = sF1i4L20;
wire sF1i5L20, cF1i5L20;
FA F1i5L20( sF1i5L20,cF1i5L20,F1i5L20_inp1,F1i5L20_inp2,F1i5L20_inp3 );

wire F1i5L21_inp1, F1i5L21_inp2, F1i5L21_inp3;
assign F1i5L21_inp1 = cF1i4L20;
assign F1i5L21_inp2 = cF2i4L20;
assign F1i5L21_inp3 = sF1i4L21;
wire sF1i5L21, cF1i5L21;
FA F1i5L21( sF1i5L21,cF1i5L21,F1i5L21_inp1,F1i5L21_inp2,F1i5L21_inp3 );

wire F1i5L22_inp1, F1i5L22_inp2, F1i5L22_inp3;
assign F1i5L22_inp1 = cF1i4L21;
assign F1i5L22_inp2 = cF2i4L21;
assign F1i5L22_inp3 = sF1i4L22;
wire sF1i5L22, cF1i5L22;
FA F1i5L22( sF1i5L22,cF1i5L22,F1i5L22_inp1,F1i5L22_inp2,F1i5L22_inp3 );

wire F1i5L23_inp1, F1i5L23_inp2, F1i5L23_inp3;
assign F1i5L23_inp1 = cF1i4L22;
assign F1i5L23_inp2 = cF2i4L22;
assign F1i5L23_inp3 = sF1i4L23;
wire sF1i5L23, cF1i5L23;
FA F1i5L23( sF1i5L23,cF1i5L23,F1i5L23_inp1,F1i5L23_inp2,F1i5L23_inp3 );

wire F1i5L24_inp1, F1i5L24_inp2, F1i5L24_inp3;
assign F1i5L24_inp1 = cF1i4L23;
assign F1i5L24_inp2 = cF2i4L23;
assign F1i5L24_inp3 = sF1i4L24;
wire sF1i5L24, cF1i5L24;
FA F1i5L24( sF1i5L24,cF1i5L24,F1i5L24_inp1,F1i5L24_inp2,F1i5L24_inp3 );

wire F1i5L25_inp1, F1i5L25_inp2, F1i5L25_inp3;
assign F1i5L25_inp1 = PP[15][10];
assign F1i5L25_inp2 = cF1i4L24;
assign F1i5L25_inp3 = cF2i4L24;
wire sF1i5L25, cF1i5L25;
FA F1i5L25( sF1i5L25,cF1i5L25,F1i5L25_inp1,F1i5L25_inp2,F1i5L25_inp3 );

wire F1i5L26_inp1, F1i5L26_inp2, F1i5L26_inp3;
assign F1i5L26_inp1 = ~PP[13][13];
assign F1i5L26_inp2 = PP[14][12];
assign F1i5L26_inp3 = PP[15][11];
wire sF1i5L26, cF1i5L26;
FA F1i5L26( sF1i5L26,cF1i5L26,F1i5L26_inp1,F1i5L26_inp2,F1i5L26_inp3 );



///////////// Iteration Number =6///////////////////





wire Hi6L2_inp1, Hi6L2_inp2;
assign Hi6L2_inp1 = PP[0][2];
assign Hi6L2_inp2 = PP[1][1];
wire sHi6L2, cHi6L2;
HA Hi6L2 ( sHi6L2,cHi6L2,Hi6L2_inp1,Hi6L2_inp2 );

wire F1i6L3_inp1, F1i6L3_inp2, F1i6L3_inp3;
assign F1i6L3_inp1 = PP[2][1];
assign F1i6L3_inp2 = PP[3][0];
assign F1i6L3_inp3 = sHi5L3;
wire sF1i6L3, cF1i6L3;
FA F1i6L3( sF1i6L3,cF1i6L3,F1i6L3_inp1,F1i6L3_inp2,F1i6L3_inp3 );

wire F1i6L4_inp1, F1i6L4_inp2, F1i6L4_inp3;
assign F1i6L4_inp1 = sHi4L4;
assign F1i6L4_inp2 = cHi5L3;
assign F1i6L4_inp3 = sF1i5L4;
wire sF1i6L4, cF1i6L4;
FA F1i6L4( sF1i6L4,cF1i6L4,F1i6L4_inp1,F1i6L4_inp2,F1i6L4_inp3 );

wire F1i6L5_inp1, F1i6L5_inp2, F1i6L5_inp3;
assign F1i6L5_inp1 = sHi4L5;
assign F1i6L5_inp2 = cF1i5L4;
assign F1i6L5_inp3 = sF1i5L5;
wire sF1i6L5, cF1i6L5;
FA F1i6L5( sF1i6L5,cF1i6L5,F1i6L5_inp1,F1i6L5_inp2,F1i6L5_inp3 );

wire F1i6L6_inp1, F1i6L6_inp2, F1i6L6_inp3;
assign F1i6L6_inp1 = sF2i4L6;
assign F1i6L6_inp2 = cF1i5L5;
assign F1i6L6_inp3 = sF1i5L6;
wire sF1i6L6, cF1i6L6;
FA F1i6L6( sF1i6L6,cF1i6L6,F1i6L6_inp1,F1i6L6_inp2,F1i6L6_inp3 );

wire F1i6L7_inp1, F1i6L7_inp2, F1i6L7_inp3;
assign F1i6L7_inp1 = sF2i4L7;
assign F1i6L7_inp2 = cF1i5L6;
assign F1i6L7_inp3 = sF1i5L7;
wire sF1i6L7, cF1i6L7;
FA F1i6L7( sF1i6L7,cF1i6L7,F1i6L7_inp1,F1i6L7_inp2,F1i6L7_inp3 );

wire F1i6L8_inp1, F1i6L8_inp2, F1i6L8_inp3;
assign F1i6L8_inp1 = sF2i4L8;
assign F1i6L8_inp2 = cF1i5L7;
assign F1i6L8_inp3 = sF1i5L8;
wire sF1i6L8, cF1i6L8;
FA F1i6L8( sF1i6L8,cF1i6L8,F1i6L8_inp1,F1i6L8_inp2,F1i6L8_inp3 );

wire F1i6L9_inp1, F1i6L9_inp2, F1i6L9_inp3;
assign F1i6L9_inp1 = sF2i4L9;
assign F1i6L9_inp2 = cF1i5L8;
assign F1i6L9_inp3 = sF1i5L9;
wire sF1i6L9, cF1i6L9;
FA F1i6L9( sF1i6L9,cF1i6L9,F1i6L9_inp1,F1i6L9_inp2,F1i6L9_inp3 );

wire F1i6L10_inp1, F1i6L10_inp2, F1i6L10_inp3;
assign F1i6L10_inp1 = sF2i4L10;
assign F1i6L10_inp2 = cF1i5L9;
assign F1i6L10_inp3 = sF1i5L10;
wire sF1i6L10, cF1i6L10;
FA F1i6L10( sF1i6L10,cF1i6L10,F1i6L10_inp1,F1i6L10_inp2,F1i6L10_inp3 );

wire F1i6L11_inp1, F1i6L11_inp2, F1i6L11_inp3;
assign F1i6L11_inp1 = sF2i4L11;
assign F1i6L11_inp2 = cF1i5L10;
assign F1i6L11_inp3 = sF1i5L11;
wire sF1i6L11, cF1i6L11;
FA F1i6L11( sF1i6L11,cF1i6L11,F1i6L11_inp1,F1i6L11_inp2,F1i6L11_inp3 );

wire F1i6L12_inp1, F1i6L12_inp2, F1i6L12_inp3;
assign F1i6L12_inp1 = sF2i4L12;
assign F1i6L12_inp2 = cF1i5L11;
assign F1i6L12_inp3 = sF1i5L12;
wire sF1i6L12, cF1i6L12;
FA F1i6L12( sF1i6L12,cF1i6L12,F1i6L12_inp1,F1i6L12_inp2,F1i6L12_inp3 );

wire F1i6L13_inp1, F1i6L13_inp2, F1i6L13_inp3;
assign F1i6L13_inp1 = sF2i4L13;
assign F1i6L13_inp2 = cF1i5L12;
assign F1i6L13_inp3 = sF1i5L13;
wire sF1i6L13, cF1i6L13;
FA F1i6L13( sF1i6L13,cF1i6L13,F1i6L13_inp1,F1i6L13_inp2,F1i6L13_inp3 );

wire F1i6L14_inp1, F1i6L14_inp2, F1i6L14_inp3;
assign F1i6L14_inp1 = sF2i4L14;
assign F1i6L14_inp2 = cF1i5L13;
assign F1i6L14_inp3 = sF1i5L14;
wire sF1i6L14, cF1i6L14;
FA F1i6L14( sF1i6L14,cF1i6L14,F1i6L14_inp1,F1i6L14_inp2,F1i6L14_inp3 );

wire F1i6L15_inp1, F1i6L15_inp2, F1i6L15_inp3;
assign F1i6L15_inp1 = sF2i4L15;
assign F1i6L15_inp2 = cF1i5L14;
assign F1i6L15_inp3 = sF1i5L15;
wire sF1i6L15, cF1i6L15;
FA F1i6L15( sF1i6L15,cF1i6L15,F1i6L15_inp1,F1i6L15_inp2,F1i6L15_inp3 );

wire F1i6L16_inp1, F1i6L16_inp2, F1i6L16_inp3;
assign F1i6L16_inp1 = sF2i4L16;
assign F1i6L16_inp2 = cF1i5L15;
assign F1i6L16_inp3 = sF1i5L16;
wire sF1i6L16, cF1i6L16;
FA F1i6L16( sF1i6L16,cF1i6L16,F1i6L16_inp1,F1i6L16_inp2,F1i6L16_inp3 );

wire F1i6L17_inp1, F1i6L17_inp2, F1i6L17_inp3;
assign F1i6L17_inp1 = sF2i4L17;
assign F1i6L17_inp2 = cF1i5L16;
assign F1i6L17_inp3 = sF1i5L17;
wire sF1i6L17, cF1i6L17;
FA F1i6L17( sF1i6L17,cF1i6L17,F1i6L17_inp1,F1i6L17_inp2,F1i6L17_inp3 );

wire F1i6L18_inp1, F1i6L18_inp2, F1i6L18_inp3;
assign F1i6L18_inp1 = sF2i4L18;
assign F1i6L18_inp2 = cF1i5L17;
assign F1i6L18_inp3 = sF1i5L18;
wire sF1i6L18, cF1i6L18;
FA F1i6L18( sF1i6L18,cF1i6L18,F1i6L18_inp1,F1i6L18_inp2,F1i6L18_inp3 );

wire F1i6L19_inp1, F1i6L19_inp2, F1i6L19_inp3;
assign F1i6L19_inp1 = sF2i4L19;
assign F1i6L19_inp2 = cF1i5L18;
assign F1i6L19_inp3 = sF1i5L19;
wire sF1i6L19, cF1i6L19;
FA F1i6L19( sF1i6L19,cF1i6L19,F1i6L19_inp1,F1i6L19_inp2,F1i6L19_inp3 );

wire F1i6L20_inp1, F1i6L20_inp2, F1i6L20_inp3;
assign F1i6L20_inp1 = sF2i4L20;
assign F1i6L20_inp2 = cF1i5L19;
assign F1i6L20_inp3 = sF1i5L20;
wire sF1i6L20, cF1i6L20;
FA F1i6L20( sF1i6L20,cF1i6L20,F1i6L20_inp1,F1i6L20_inp2,F1i6L20_inp3 );

wire F1i6L21_inp1, F1i6L21_inp2, F1i6L21_inp3;
assign F1i6L21_inp1 = sF2i4L21;
assign F1i6L21_inp2 = cF1i5L20;
assign F1i6L21_inp3 = sF1i5L21;
wire sF1i6L21, cF1i6L21;
FA F1i6L21( sF1i6L21,cF1i6L21,F1i6L21_inp1,F1i6L21_inp2,F1i6L21_inp3 );

wire F1i6L22_inp1, F1i6L22_inp2, F1i6L22_inp3;
assign F1i6L22_inp1 = sF2i4L22;
assign F1i6L22_inp2 = cF1i5L21;
assign F1i6L22_inp3 = sF1i5L22;
wire sF1i6L22, cF1i6L22;
FA F1i6L22( sF1i6L22,cF1i6L22,F1i6L22_inp1,F1i6L22_inp2,F1i6L22_inp3 );

wire F1i6L23_inp1, F1i6L23_inp2, F1i6L23_inp3;
assign F1i6L23_inp1 = sF2i4L23;
assign F1i6L23_inp2 = cF1i5L22;
assign F1i6L23_inp3 = sF1i5L23;
wire sF1i6L23, cF1i6L23;
FA F1i6L23( sF1i6L23,cF1i6L23,F1i6L23_inp1,F1i6L23_inp2,F1i6L23_inp3 );

wire F1i6L24_inp1, F1i6L24_inp2, F1i6L24_inp3;
assign F1i6L24_inp1 = sF2i4L24;
assign F1i6L24_inp2 = cF1i5L23;
assign F1i6L24_inp3 = sF1i5L24;
wire sF1i6L24, cF1i6L24;
FA F1i6L24( sF1i6L24,cF1i6L24,F1i6L24_inp1,F1i6L24_inp2,F1i6L24_inp3 );

wire F1i6L25_inp1, F1i6L25_inp2, F1i6L25_inp3;
assign F1i6L25_inp1 = sF1i4L25;
assign F1i6L25_inp2 = cF1i5L24;
assign F1i6L25_inp3 = sF1i5L25;
wire sF1i6L25, cF1i6L25;
FA F1i6L25( sF1i6L25,cF1i6L25,F1i6L25_inp1,F1i6L25_inp2,F1i6L25_inp3 );

wire F1i6L26_inp1, F1i6L26_inp2, F1i6L26_inp3;
assign F1i6L26_inp1 = cF1i4L25;
assign F1i6L26_inp2 = cF1i5L25;
assign F1i6L26_inp3 = sF1i5L26;
wire sF1i6L26, cF1i6L26;
FA F1i6L26( sF1i6L26,cF1i6L26,F1i6L26_inp1,F1i6L26_inp2,F1i6L26_inp3 );

wire F1i6L27_inp1, F1i6L27_inp2, F1i6L27_inp3;
assign F1i6L27_inp1 = ~PP[14][13];
assign F1i6L27_inp2 = PP[15][12];
assign F1i6L27_inp3 = cF1i5L26;
wire sF1i6L27, cF1i6L27;
FA F1i6L27( sF1i6L27,cF1i6L27,F1i6L27_inp1,F1i6L27_inp2,F1i6L27_inp3 );


assign out1 ={{CV[29]},{~PP[15][13]},{cF1i6L26},{cF1i6L25},{cF1i6L24},{cF1i6L23},{cF1i6L22},{cF1i6L21},{cF1i6L20},{cF1i6L19},{cF1i6L18},{cF1i6L17},{cF1i6L16},{cF1i6L15},{cF1i6L14},{cF1i6L13},{cF1i6L12},{cF1i6L11},{cF1i6L10},{cF1i6L9},{cF1i6L8},{cF1i6L7},{cF1i6L6},{cF1i6L5},{cF1i6L4},{cF1i6L3},{cHi6L2},{PP[2][0]},{PP[0][1]},{PP[0][0]}};
assign out2 ={{1'b0},{cF1i6L27},{sF1i6L27},{sF1i6L26},{sF1i6L25},{sF1i6L24},{sF1i6L23},{sF1i6L22},{sF1i6L21},{sF1i6L20},{sF1i6L19},{sF1i6L18},{sF1i6L17},{sF1i6L16},{sF1i6L15},{sF1i6L14},{sF1i6L13},{sF1i6L12},{sF1i6L11},{sF1i6L10},{sF1i6L9},{sF1i6L8},{sF1i6L7},{sF1i6L6},{sF1i6L5},{sF1i6L4},{sF1i6L3},{sHi6L2},{PP[1][0]},{1'b0}} ;
endmodule